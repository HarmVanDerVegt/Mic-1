library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

entity control_store is

  port (
    address     : in  std_logic_vector(8 downto 0);
    test        : out std_logic_vector(35 downto 0);
    instruction : out std_logic_vector(35 downto 0));

end entity control_store;

architecture control_store_ar of control_store is
  component decoder is
    generic (
      input_count  : natural := 9;
      output_count : natural := 512);
    port (
      input  : in  std_logic_vector(input_count - 1 downto 0);
      output : out std_logic_vector(output_count - 1 downto 0));
  end component decoder;

  component rom is
    generic (
      bits  : natural;
      value : std_logic_vector(36 -1 downto 0));
    port (
      enable_o : in  std_logic;
      output   : out std_logic_vector(bits -1 downto 0));
  end component rom;

  signal mem_enable_lines : std_logic_vector(511 downto 0);
  type mem_array_type is array (35 downto 0) of std_logic_vector(511 downto 0);
  signal mem_array        : mem_array_type;
  signal temp_instruction : std_logic_vector(35 downto 0) := (others => '0');

begin  -- architecture control_store_ar

  decoder1 : entity work.decoder
    generic map (
      input_count  => 9,
      output_count => 512)
    port map (
      input  => address,
      output => mem_enable_lines);

  rom0 : entity work.rom
    generic map (
      bits  => 36,
      value => "000100100011010001010110011110000000")
    port map (
      enable_o   => mem_enable_lines(0),
      output(0)  => mem_array(0)(0),
      output(1)  => mem_array(1)(0),
      output(2)  => mem_array(2)(0),
      output(3)  => mem_array(3)(0),
      output(4)  => mem_array(4)(0),
      output(5)  => mem_array(5)(0),
      output(6)  => mem_array(6)(0),
      output(7)  => mem_array(7)(0),
      output(8)  => mem_array(8)(0),
      output(9)  => mem_array(9)(0),
      output(10) => mem_array(10)(0),
      output(11) => mem_array(11)(0),
      output(12) => mem_array(12)(0),
      output(13) => mem_array(13)(0),
      output(14) => mem_array(14)(0),
      output(15) => mem_array(15)(0),
      output(16) => mem_array(16)(0),
      output(17) => mem_array(17)(0),
      output(18) => mem_array(18)(0),
      output(19) => mem_array(19)(0),
      output(20) => mem_array(20)(0),
      output(21) => mem_array(21)(0),
      output(22) => mem_array(22)(0),
      output(23) => mem_array(23)(0),
      output(24) => mem_array(24)(0),
      output(25) => mem_array(25)(0),
      output(26) => mem_array(26)(0),
      output(27) => mem_array(27)(0),
      output(28) => mem_array(28)(0),
      output(29) => mem_array(29)(0),
      output(30) => mem_array(30)(0),
      output(31) => mem_array(31)(0),
      output(32) => mem_array(32)(0),
      output(33) => mem_array(33)(0),
      output(34) => mem_array(34)(0),
      output(35) => mem_array(35)(0)
      );
  rom1 : entity work.rom
    generic map (
      bits  => 36,
      value => "000100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(1),
      output(0)  => mem_array(0)(1),
      output(1)  => mem_array(1)(1),
      output(2)  => mem_array(2)(1),
      output(3)  => mem_array(3)(1),
      output(4)  => mem_array(4)(1),
      output(5)  => mem_array(5)(1),
      output(6)  => mem_array(6)(1),
      output(7)  => mem_array(7)(1),
      output(8)  => mem_array(8)(1),
      output(9)  => mem_array(9)(1),
      output(10) => mem_array(10)(1),
      output(11) => mem_array(11)(1),
      output(12) => mem_array(12)(1),
      output(13) => mem_array(13)(1),
      output(14) => mem_array(14)(1),
      output(15) => mem_array(15)(1),
      output(16) => mem_array(16)(1),
      output(17) => mem_array(17)(1),
      output(18) => mem_array(18)(1),
      output(19) => mem_array(19)(1),
      output(20) => mem_array(20)(1),
      output(21) => mem_array(21)(1),
      output(22) => mem_array(22)(1),
      output(23) => mem_array(23)(1),
      output(24) => mem_array(24)(1),
      output(25) => mem_array(25)(1),
      output(26) => mem_array(26)(1),
      output(27) => mem_array(27)(1),
      output(28) => mem_array(28)(1),
      output(29) => mem_array(29)(1),
      output(30) => mem_array(30)(1),
      output(31) => mem_array(31)(1),
      output(32) => mem_array(32)(1),
      output(33) => mem_array(33)(1),
      output(34) => mem_array(34)(1),
      output(35) => mem_array(35)(1)
      );
  rom2 : entity work.rom
    generic map (
      bits  => 36,
      value => "001000000000001101010000001000000001")
    port map (
      enable_o   => mem_enable_lines(2),
      output(0)  => mem_array(0)(2),
      output(1)  => mem_array(1)(2),
      output(2)  => mem_array(2)(2),
      output(3)  => mem_array(3)(2),
      output(4)  => mem_array(4)(2),
      output(5)  => mem_array(5)(2),
      output(6)  => mem_array(6)(2),
      output(7)  => mem_array(7)(2),
      output(8)  => mem_array(8)(2),
      output(9)  => mem_array(9)(2),
      output(10) => mem_array(10)(2),
      output(11) => mem_array(11)(2),
      output(12) => mem_array(12)(2),
      output(13) => mem_array(13)(2),
      output(14) => mem_array(14)(2),
      output(15) => mem_array(15)(2),
      output(16) => mem_array(16)(2),
      output(17) => mem_array(17)(2),
      output(18) => mem_array(18)(2),
      output(19) => mem_array(19)(2),
      output(20) => mem_array(20)(2),
      output(21) => mem_array(21)(2),
      output(22) => mem_array(22)(2),
      output(23) => mem_array(23)(2),
      output(24) => mem_array(24)(2),
      output(25) => mem_array(25)(2),
      output(26) => mem_array(26)(2),
      output(27) => mem_array(27)(2),
      output(28) => mem_array(28)(2),
      output(29) => mem_array(29)(2),
      output(30) => mem_array(30)(2),
      output(31) => mem_array(31)(2),
      output(32) => mem_array(32)(2),
      output(33) => mem_array(33)(2),
      output(34) => mem_array(34)(2),
      output(35) => mem_array(35)(2)
      );
  rom3 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000010000110101000000100001")
    port map (
      enable_o   => mem_enable_lines(3),
      output(0)  => mem_array(0)(3),
      output(1)  => mem_array(1)(3),
      output(2)  => mem_array(2)(3),
      output(3)  => mem_array(3)(3),
      output(4)  => mem_array(4)(3),
      output(5)  => mem_array(5)(3),
      output(6)  => mem_array(6)(3),
      output(7)  => mem_array(7)(3),
      output(8)  => mem_array(8)(3),
      output(9)  => mem_array(9)(3),
      output(10) => mem_array(10)(3),
      output(11) => mem_array(11)(3),
      output(12) => mem_array(12)(3),
      output(13) => mem_array(13)(3),
      output(14) => mem_array(14)(3),
      output(15) => mem_array(15)(3),
      output(16) => mem_array(16)(3),
      output(17) => mem_array(17)(3),
      output(18) => mem_array(18)(3),
      output(19) => mem_array(19)(3),
      output(20) => mem_array(20)(3),
      output(21) => mem_array(21)(3),
      output(22) => mem_array(22)(3),
      output(23) => mem_array(23)(3),
      output(24) => mem_array(24)(3),
      output(25) => mem_array(25)(3),
      output(26) => mem_array(26)(3),
      output(27) => mem_array(27)(3),
      output(28) => mem_array(28)(3),
      output(29) => mem_array(29)(3),
      output(30) => mem_array(30)(3),
      output(31) => mem_array(31)(3),
      output(32) => mem_array(32)(3),
      output(33) => mem_array(33)(3),
      output(34) => mem_array(34)(3),
      output(35) => mem_array(35)(3)
      );
  rom4 : entity work.rom
    generic map (
      bits  => 36,
      value => "000100000000001000000001010010000000")
    port map (
      enable_o   => mem_enable_lines(4),
      output(0)  => mem_array(0)(4),
      output(1)  => mem_array(1)(4),
      output(2)  => mem_array(2)(4),
      output(3)  => mem_array(3)(4),
      output(4)  => mem_array(4)(4),
      output(5)  => mem_array(5)(4),
      output(6)  => mem_array(6)(4),
      output(7)  => mem_array(7)(4),
      output(8)  => mem_array(8)(4),
      output(9)  => mem_array(9)(4),
      output(10) => mem_array(10)(4),
      output(11) => mem_array(11)(4),
      output(12) => mem_array(12)(4),
      output(13) => mem_array(13)(4),
      output(14) => mem_array(14)(4),
      output(15) => mem_array(15)(4),
      output(16) => mem_array(16)(4),
      output(17) => mem_array(17)(4),
      output(18) => mem_array(18)(4),
      output(19) => mem_array(19)(4),
      output(20) => mem_array(20)(4),
      output(21) => mem_array(21)(4),
      output(22) => mem_array(22)(4),
      output(23) => mem_array(23)(4),
      output(24) => mem_array(24)(4),
      output(25) => mem_array(25)(4),
      output(26) => mem_array(26)(4),
      output(27) => mem_array(27)(4),
      output(28) => mem_array(28)(4),
      output(29) => mem_array(29)(4),
      output(30) => mem_array(30)(4),
      output(31) => mem_array(31)(4),
      output(32) => mem_array(32)(4),
      output(33) => mem_array(33)(4),
      output(34) => mem_array(34)(4),
      output(35) => mem_array(35)(4)
      );
  rom5 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001110000000000010000001111000010")
    port map (
      enable_o   => mem_enable_lines(5),
      output(0)  => mem_array(0)(5),
      output(1)  => mem_array(1)(5),
      output(2)  => mem_array(2)(5),
      output(3)  => mem_array(3)(5),
      output(4)  => mem_array(4)(5),
      output(5)  => mem_array(5)(5),
      output(6)  => mem_array(6)(5),
      output(7)  => mem_array(7)(5),
      output(8)  => mem_array(8)(5),
      output(9)  => mem_array(9)(5),
      output(10) => mem_array(10)(5),
      output(11) => mem_array(11)(5),
      output(12) => mem_array(12)(5),
      output(13) => mem_array(13)(5),
      output(14) => mem_array(14)(5),
      output(15) => mem_array(15)(5),
      output(16) => mem_array(16)(5),
      output(17) => mem_array(17)(5),
      output(18) => mem_array(18)(5),
      output(19) => mem_array(19)(5),
      output(20) => mem_array(20)(5),
      output(21) => mem_array(21)(5),
      output(22) => mem_array(22)(5),
      output(23) => mem_array(23)(5),
      output(24) => mem_array(24)(5),
      output(25) => mem_array(25)(5),
      output(26) => mem_array(26)(5),
      output(27) => mem_array(27)(5),
      output(28) => mem_array(28)(5),
      output(29) => mem_array(29)(5),
      output(30) => mem_array(30)(5),
      output(31) => mem_array(31)(5),
      output(32) => mem_array(32)(5),
      output(33) => mem_array(33)(5),
      output(34) => mem_array(34)(5),
      output(35) => mem_array(35)(5)
      );
  rom6 : entity work.rom
    generic map (
      bits  => 36,
      value => "000101000000000000000011000000010100")
    port map (
      enable_o   => mem_enable_lines(6),
      output(0)  => mem_array(0)(6),
      output(1)  => mem_array(1)(6),
      output(2)  => mem_array(2)(6),
      output(3)  => mem_array(3)(6),
      output(4)  => mem_array(4)(6),
      output(5)  => mem_array(5)(6),
      output(6)  => mem_array(6)(6),
      output(7)  => mem_array(7)(6),
      output(8)  => mem_array(8)(6),
      output(9)  => mem_array(9)(6),
      output(10) => mem_array(10)(6),
      output(11) => mem_array(11)(6),
      output(12) => mem_array(12)(6),
      output(13) => mem_array(13)(6),
      output(14) => mem_array(14)(6),
      output(15) => mem_array(15)(6),
      output(16) => mem_array(16)(6),
      output(17) => mem_array(17)(6),
      output(18) => mem_array(18)(6),
      output(19) => mem_array(19)(6),
      output(20) => mem_array(20)(6),
      output(21) => mem_array(21)(6),
      output(22) => mem_array(22)(6),
      output(23) => mem_array(23)(6),
      output(24) => mem_array(24)(6),
      output(25) => mem_array(25)(6),
      output(26) => mem_array(26)(6),
      output(27) => mem_array(27)(6),
      output(28) => mem_array(28)(6),
      output(29) => mem_array(29)(6),
      output(30) => mem_array(30)(6),
      output(31) => mem_array(31)(6),
      output(32) => mem_array(32)(6),
      output(33) => mem_array(33)(6),
      output(34) => mem_array(34)(6),
      output(35) => mem_array(35)(6)
      );
  rom7 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000000000011100000000000100000011")
    port map (
      enable_o   => mem_enable_lines(7),
      output(0)  => mem_array(0)(7),
      output(1)  => mem_array(1)(7),
      output(2)  => mem_array(2)(7),
      output(3)  => mem_array(3)(7),
      output(4)  => mem_array(4)(7),
      output(5)  => mem_array(5)(7),
      output(6)  => mem_array(6)(7),
      output(7)  => mem_array(7)(7),
      output(8)  => mem_array(8)(7),
      output(9)  => mem_array(9)(7),
      output(10) => mem_array(10)(7),
      output(11) => mem_array(11)(7),
      output(12) => mem_array(12)(7),
      output(13) => mem_array(13)(7),
      output(14) => mem_array(14)(7),
      output(15) => mem_array(15)(7),
      output(16) => mem_array(16)(7),
      output(17) => mem_array(17)(7),
      output(18) => mem_array(18)(7),
      output(19) => mem_array(19)(7),
      output(20) => mem_array(20)(7),
      output(21) => mem_array(21)(7),
      output(22) => mem_array(22)(7),
      output(23) => mem_array(23)(7),
      output(24) => mem_array(24)(7),
      output(25) => mem_array(25)(7),
      output(26) => mem_array(26)(7),
      output(27) => mem_array(27)(7),
      output(28) => mem_array(28)(7),
      output(29) => mem_array(29)(7),
      output(30) => mem_array(30)(7),
      output(31) => mem_array(31)(7),
      output(32) => mem_array(32)(7),
      output(33) => mem_array(33)(7),
      output(34) => mem_array(34)(7),
      output(35) => mem_array(35)(7)
      );
  rom8 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100100001010000000000000001000000")
    port map (
      enable_o   => mem_enable_lines(8),
      output(0)  => mem_array(0)(8),
      output(1)  => mem_array(1)(8),
      output(2)  => mem_array(2)(8),
      output(3)  => mem_array(3)(8),
      output(4)  => mem_array(4)(8),
      output(5)  => mem_array(5)(8),
      output(6)  => mem_array(6)(8),
      output(7)  => mem_array(7)(8),
      output(8)  => mem_array(8)(8),
      output(9)  => mem_array(9)(8),
      output(10) => mem_array(10)(8),
      output(11) => mem_array(11)(8),
      output(12) => mem_array(12)(8),
      output(13) => mem_array(13)(8),
      output(14) => mem_array(14)(8),
      output(15) => mem_array(15)(8),
      output(16) => mem_array(16)(8),
      output(17) => mem_array(17)(8),
      output(18) => mem_array(18)(8),
      output(19) => mem_array(19)(8),
      output(20) => mem_array(20)(8),
      output(21) => mem_array(21)(8),
      output(22) => mem_array(22)(8),
      output(23) => mem_array(23)(8),
      output(24) => mem_array(24)(8),
      output(25) => mem_array(25)(8),
      output(26) => mem_array(26)(8),
      output(27) => mem_array(27)(8),
      output(28) => mem_array(28)(8),
      output(29) => mem_array(29)(8),
      output(30) => mem_array(30)(8),
      output(31) => mem_array(31)(8),
      output(32) => mem_array(32)(8),
      output(33) => mem_array(33)(8),
      output(34) => mem_array(34)(8),
      output(35) => mem_array(35)(8)
      );
  rom9 : entity work.rom
    generic map (
      bits  => 36,
      value => "000101001000000000000111000000000001")
    port map (
      enable_o   => mem_enable_lines(9),
      output(0)  => mem_array(0)(9),
      output(1)  => mem_array(1)(9),
      output(2)  => mem_array(2)(9),
      output(3)  => mem_array(3)(9),
      output(4)  => mem_array(4)(9),
      output(5)  => mem_array(5)(9),
      output(6)  => mem_array(6)(9),
      output(7)  => mem_array(7)(9),
      output(8)  => mem_array(8)(9),
      output(9)  => mem_array(9)(9),
      output(10) => mem_array(10)(9),
      output(11) => mem_array(11)(9),
      output(12) => mem_array(12)(9),
      output(13) => mem_array(13)(9),
      output(14) => mem_array(14)(9),
      output(15) => mem_array(15)(9),
      output(16) => mem_array(16)(9),
      output(17) => mem_array(17)(9),
      output(18) => mem_array(18)(9),
      output(19) => mem_array(19)(9),
      output(20) => mem_array(20)(9),
      output(21) => mem_array(21)(9),
      output(22) => mem_array(22)(9),
      output(23) => mem_array(23)(9),
      output(24) => mem_array(24)(9),
      output(25) => mem_array(25)(9),
      output(26) => mem_array(26)(9),
      output(27) => mem_array(27)(9),
      output(28) => mem_array(28)(9),
      output(29) => mem_array(29)(9),
      output(30) => mem_array(30)(9),
      output(31) => mem_array(31)(9),
      output(32) => mem_array(32)(9),
      output(33) => mem_array(33)(9),
      output(34) => mem_array(34)(9),
      output(35) => mem_array(35)(9)
      );
  rom10 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001100001000010100000000000000")
    port map (
      enable_o   => mem_enable_lines(10),
      output(0)  => mem_array(0)(10),
      output(1)  => mem_array(1)(10),
      output(2)  => mem_array(2)(10),
      output(3)  => mem_array(3)(10),
      output(4)  => mem_array(4)(10),
      output(5)  => mem_array(5)(10),
      output(6)  => mem_array(6)(10),
      output(7)  => mem_array(7)(10),
      output(8)  => mem_array(8)(10),
      output(9)  => mem_array(9)(10),
      output(10) => mem_array(10)(10),
      output(11) => mem_array(11)(10),
      output(12) => mem_array(12)(10),
      output(13) => mem_array(13)(10),
      output(14) => mem_array(14)(10),
      output(15) => mem_array(15)(10),
      output(16) => mem_array(16)(10),
      output(17) => mem_array(17)(10),
      output(18) => mem_array(18)(10),
      output(19) => mem_array(19)(10),
      output(20) => mem_array(20)(10),
      output(21) => mem_array(21)(10),
      output(22) => mem_array(22)(10),
      output(23) => mem_array(23)(10),
      output(24) => mem_array(24)(10),
      output(25) => mem_array(25)(10),
      output(26) => mem_array(26)(10),
      output(27) => mem_array(27)(10),
      output(28) => mem_array(28)(10),
      output(29) => mem_array(29)(10),
      output(30) => mem_array(30)(10),
      output(31) => mem_array(31)(10),
      output(32) => mem_array(32)(10),
      output(33) => mem_array(33)(10),
      output(34) => mem_array(34)(10),
      output(35) => mem_array(35)(10)
      );
  rom11 : entity work.rom
    generic map (
      bits  => 36,
      value => "010100000001010010000000000001110000")
    port map (
      enable_o   => mem_enable_lines(11),
      output(0)  => mem_array(0)(11),
      output(1)  => mem_array(1)(11),
      output(2)  => mem_array(2)(11),
      output(3)  => mem_array(3)(11),
      output(4)  => mem_array(4)(11),
      output(5)  => mem_array(5)(11),
      output(6)  => mem_array(6)(11),
      output(7)  => mem_array(7)(11),
      output(8)  => mem_array(8)(11),
      output(9)  => mem_array(9)(11),
      output(10) => mem_array(10)(11),
      output(11) => mem_array(11)(11),
      output(12) => mem_array(12)(11),
      output(13) => mem_array(13)(11),
      output(14) => mem_array(14)(11),
      output(15) => mem_array(15)(11),
      output(16) => mem_array(16)(11),
      output(17) => mem_array(17)(11),
      output(18) => mem_array(18)(11),
      output(19) => mem_array(19)(11),
      output(20) => mem_array(20)(11),
      output(21) => mem_array(21)(11),
      output(22) => mem_array(22)(11),
      output(23) => mem_array(23)(11),
      output(24) => mem_array(24)(11),
      output(25) => mem_array(25)(11),
      output(26) => mem_array(26)(11),
      output(27) => mem_array(27)(11),
      output(28) => mem_array(28)(11),
      output(29) => mem_array(29)(11),
      output(30) => mem_array(30)(11),
      output(31) => mem_array(31)(11),
      output(32) => mem_array(32)(11),
      output(33) => mem_array(33)(11),
      output(34) => mem_array(34)(11),
      output(35) => mem_array(35)(11)
      );
  rom12 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000010000000111000010000101000000")
    port map (
      enable_o   => mem_enable_lines(12),
      output(0)  => mem_array(0)(12),
      output(1)  => mem_array(1)(12),
      output(2)  => mem_array(2)(12),
      output(3)  => mem_array(3)(12),
      output(4)  => mem_array(4)(12),
      output(5)  => mem_array(5)(12),
      output(6)  => mem_array(6)(12),
      output(7)  => mem_array(7)(12),
      output(8)  => mem_array(8)(12),
      output(9)  => mem_array(9)(12),
      output(10) => mem_array(10)(12),
      output(11) => mem_array(11)(12),
      output(12) => mem_array(12)(12),
      output(13) => mem_array(13)(12),
      output(14) => mem_array(14)(12),
      output(15) => mem_array(15)(12),
      output(16) => mem_array(16)(12),
      output(17) => mem_array(17)(12),
      output(18) => mem_array(18)(12),
      output(19) => mem_array(19)(12),
      output(20) => mem_array(20)(12),
      output(21) => mem_array(21)(12),
      output(22) => mem_array(22)(12),
      output(23) => mem_array(23)(12),
      output(24) => mem_array(24)(12),
      output(25) => mem_array(25)(12),
      output(26) => mem_array(26)(12),
      output(27) => mem_array(27)(12),
      output(28) => mem_array(28)(12),
      output(29) => mem_array(29)(12),
      output(30) => mem_array(30)(12),
      output(31) => mem_array(31)(12),
      output(32) => mem_array(32)(12),
      output(33) => mem_array(33)(12),
      output(34) => mem_array(34)(12),
      output(35) => mem_array(35)(12)
      );
  rom13 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000001000000010100000000010100")
    port map (
      enable_o   => mem_enable_lines(13),
      output(0)  => mem_array(0)(13),
      output(1)  => mem_array(1)(13),
      output(2)  => mem_array(2)(13),
      output(3)  => mem_array(3)(13),
      output(4)  => mem_array(4)(13),
      output(5)  => mem_array(5)(13),
      output(6)  => mem_array(6)(13),
      output(7)  => mem_array(7)(13),
      output(8)  => mem_array(8)(13),
      output(9)  => mem_array(9)(13),
      output(10) => mem_array(10)(13),
      output(11) => mem_array(11)(13),
      output(12) => mem_array(12)(13),
      output(13) => mem_array(13)(13),
      output(14) => mem_array(14)(13),
      output(15) => mem_array(15)(13),
      output(16) => mem_array(16)(13),
      output(17) => mem_array(17)(13),
      output(18) => mem_array(18)(13),
      output(19) => mem_array(19)(13),
      output(20) => mem_array(20)(13),
      output(21) => mem_array(21)(13),
      output(22) => mem_array(22)(13),
      output(23) => mem_array(23)(13),
      output(24) => mem_array(24)(13),
      output(25) => mem_array(25)(13),
      output(26) => mem_array(26)(13),
      output(27) => mem_array(27)(13),
      output(28) => mem_array(28)(13),
      output(29) => mem_array(29)(13),
      output(30) => mem_array(30)(13),
      output(31) => mem_array(31)(13),
      output(32) => mem_array(32)(13),
      output(33) => mem_array(33)(13),
      output(34) => mem_array(34)(13),
      output(35) => mem_array(35)(13)
      );
  rom14 : entity work.rom
    generic map (
      bits  => 36,
      value => "011100000000011010000000000000000000")
    port map (
      enable_o   => mem_enable_lines(14),
      output(0)  => mem_array(0)(14),
      output(1)  => mem_array(1)(14),
      output(2)  => mem_array(2)(14),
      output(3)  => mem_array(3)(14),
      output(4)  => mem_array(4)(14),
      output(5)  => mem_array(5)(14),
      output(6)  => mem_array(6)(14),
      output(7)  => mem_array(7)(14),
      output(8)  => mem_array(8)(14),
      output(9)  => mem_array(9)(14),
      output(10) => mem_array(10)(14),
      output(11) => mem_array(11)(14),
      output(12) => mem_array(12)(14),
      output(13) => mem_array(13)(14),
      output(14) => mem_array(14)(14),
      output(15) => mem_array(15)(14),
      output(16) => mem_array(16)(14),
      output(17) => mem_array(17)(14),
      output(18) => mem_array(18)(14),
      output(19) => mem_array(19)(14),
      output(20) => mem_array(20)(14),
      output(21) => mem_array(21)(14),
      output(22) => mem_array(22)(14),
      output(23) => mem_array(23)(14),
      output(24) => mem_array(24)(14),
      output(25) => mem_array(25)(14),
      output(26) => mem_array(26)(14),
      output(27) => mem_array(27)(14),
      output(28) => mem_array(28)(14),
      output(29) => mem_array(29)(14),
      output(30) => mem_array(30)(14),
      output(31) => mem_array(31)(14),
      output(32) => mem_array(32)(14),
      output(33) => mem_array(33)(14),
      output(34) => mem_array(34)(14),
      output(35) => mem_array(35)(14)
      );
  rom15 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000010000000101000010")
    port map (
      enable_o   => mem_enable_lines(15),
      output(0)  => mem_array(0)(15),
      output(1)  => mem_array(1)(15),
      output(2)  => mem_array(2)(15),
      output(3)  => mem_array(3)(15),
      output(4)  => mem_array(4)(15),
      output(5)  => mem_array(5)(15),
      output(6)  => mem_array(6)(15),
      output(7)  => mem_array(7)(15),
      output(8)  => mem_array(8)(15),
      output(9)  => mem_array(9)(15),
      output(10) => mem_array(10)(15),
      output(11) => mem_array(11)(15),
      output(12) => mem_array(12)(15),
      output(13) => mem_array(13)(15),
      output(14) => mem_array(14)(15),
      output(15) => mem_array(15)(15),
      output(16) => mem_array(16)(15),
      output(17) => mem_array(17)(15),
      output(18) => mem_array(18)(15),
      output(19) => mem_array(19)(15),
      output(20) => mem_array(20)(15),
      output(21) => mem_array(21)(15),
      output(22) => mem_array(22)(15),
      output(23) => mem_array(23)(15),
      output(24) => mem_array(24)(15),
      output(25) => mem_array(25)(15),
      output(26) => mem_array(26)(15),
      output(27) => mem_array(27)(15),
      output(28) => mem_array(28)(15),
      output(29) => mem_array(29)(15),
      output(30) => mem_array(30)(15),
      output(31) => mem_array(31)(15),
      output(32) => mem_array(32)(15),
      output(33) => mem_array(33)(15),
      output(34) => mem_array(34)(15),
      output(35) => mem_array(35)(15)
      );
  rom16 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111100000010100")
    port map (
      enable_o   => mem_enable_lines(16),
      output(0)  => mem_array(0)(16),
      output(1)  => mem_array(1)(16),
      output(2)  => mem_array(2)(16),
      output(3)  => mem_array(3)(16),
      output(4)  => mem_array(4)(16),
      output(5)  => mem_array(5)(16),
      output(6)  => mem_array(6)(16),
      output(7)  => mem_array(7)(16),
      output(8)  => mem_array(8)(16),
      output(9)  => mem_array(9)(16),
      output(10) => mem_array(10)(16),
      output(11) => mem_array(11)(16),
      output(12) => mem_array(12)(16),
      output(13) => mem_array(13)(16),
      output(14) => mem_array(14)(16),
      output(15) => mem_array(15)(16),
      output(16) => mem_array(16)(16),
      output(17) => mem_array(17)(16),
      output(18) => mem_array(18)(16),
      output(19) => mem_array(19)(16),
      output(20) => mem_array(20)(16),
      output(21) => mem_array(21)(16),
      output(22) => mem_array(22)(16),
      output(23) => mem_array(23)(16),
      output(24) => mem_array(24)(16),
      output(25) => mem_array(25)(16),
      output(26) => mem_array(26)(16),
      output(27) => mem_array(27)(16),
      output(28) => mem_array(28)(16),
      output(29) => mem_array(29)(16),
      output(30) => mem_array(30)(16),
      output(31) => mem_array(31)(16),
      output(32) => mem_array(32)(16),
      output(33) => mem_array(33)(16),
      output(34) => mem_array(34)(16),
      output(35) => mem_array(35)(16)
      );
  rom17 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001000010000000000100010000001")
    port map (
      enable_o   => mem_enable_lines(17),
      output(0)  => mem_array(0)(17),
      output(1)  => mem_array(1)(17),
      output(2)  => mem_array(2)(17),
      output(3)  => mem_array(3)(17),
      output(4)  => mem_array(4)(17),
      output(5)  => mem_array(5)(17),
      output(6)  => mem_array(6)(17),
      output(7)  => mem_array(7)(17),
      output(8)  => mem_array(8)(17),
      output(9)  => mem_array(9)(17),
      output(10) => mem_array(10)(17),
      output(11) => mem_array(11)(17),
      output(12) => mem_array(12)(17),
      output(13) => mem_array(13)(17),
      output(14) => mem_array(14)(17),
      output(15) => mem_array(15)(17),
      output(16) => mem_array(16)(17),
      output(17) => mem_array(17)(17),
      output(18) => mem_array(18)(17),
      output(19) => mem_array(19)(17),
      output(20) => mem_array(20)(17),
      output(21) => mem_array(21)(17),
      output(22) => mem_array(22)(17),
      output(23) => mem_array(23)(17),
      output(24) => mem_array(24)(17),
      output(25) => mem_array(25)(17),
      output(26) => mem_array(26)(17),
      output(27) => mem_array(27)(17),
      output(28) => mem_array(28)(17),
      output(29) => mem_array(29)(17),
      output(30) => mem_array(30)(17),
      output(31) => mem_array(31)(17),
      output(32) => mem_array(32)(17),
      output(33) => mem_array(33)(17),
      output(34) => mem_array(34)(17),
      output(35) => mem_array(35)(17)
      );
  rom18 : entity work.rom
    generic map (
      bits  => 36,
      value => "010010000000010000000000000010110000")
    port map (
      enable_o   => mem_enable_lines(18),
      output(0)  => mem_array(0)(18),
      output(1)  => mem_array(1)(18),
      output(2)  => mem_array(2)(18),
      output(3)  => mem_array(3)(18),
      output(4)  => mem_array(4)(18),
      output(5)  => mem_array(5)(18),
      output(6)  => mem_array(6)(18),
      output(7)  => mem_array(7)(18),
      output(8)  => mem_array(8)(18),
      output(9)  => mem_array(9)(18),
      output(10) => mem_array(10)(18),
      output(11) => mem_array(11)(18),
      output(12) => mem_array(12)(18),
      output(13) => mem_array(13)(18),
      output(14) => mem_array(14)(18),
      output(15) => mem_array(15)(18),
      output(16) => mem_array(16)(18),
      output(17) => mem_array(17)(18),
      output(18) => mem_array(18)(18),
      output(19) => mem_array(19)(18),
      output(20) => mem_array(20)(18),
      output(21) => mem_array(21)(18),
      output(22) => mem_array(22)(18),
      output(23) => mem_array(23)(18),
      output(24) => mem_array(24)(18),
      output(25) => mem_array(25)(18),
      output(26) => mem_array(26)(18),
      output(27) => mem_array(27)(18),
      output(28) => mem_array(28)(18),
      output(29) => mem_array(29)(18),
      output(30) => mem_array(30)(18),
      output(31) => mem_array(31)(18),
      output(32) => mem_array(32)(18),
      output(33) => mem_array(33)(18),
      output(34) => mem_array(34)(18),
      output(35) => mem_array(35)(18)
      );
  rom19 : entity work.rom
    generic map (
      bits  => 36,
      value => "001101010000010010000100000000001001")
    port map (
      enable_o   => mem_enable_lines(19),
      output(0)  => mem_array(0)(19),
      output(1)  => mem_array(1)(19),
      output(2)  => mem_array(2)(19),
      output(3)  => mem_array(3)(19),
      output(4)  => mem_array(4)(19),
      output(5)  => mem_array(5)(19),
      output(6)  => mem_array(6)(19),
      output(7)  => mem_array(7)(19),
      output(8)  => mem_array(8)(19),
      output(9)  => mem_array(9)(19),
      output(10) => mem_array(10)(19),
      output(11) => mem_array(11)(19),
      output(12) => mem_array(12)(19),
      output(13) => mem_array(13)(19),
      output(14) => mem_array(14)(19),
      output(15) => mem_array(15)(19),
      output(16) => mem_array(16)(19),
      output(17) => mem_array(17)(19),
      output(18) => mem_array(18)(19),
      output(19) => mem_array(19)(19),
      output(20) => mem_array(20)(19),
      output(21) => mem_array(21)(19),
      output(22) => mem_array(22)(19),
      output(23) => mem_array(23)(19),
      output(24) => mem_array(24)(19),
      output(25) => mem_array(25)(19),
      output(26) => mem_array(26)(19),
      output(27) => mem_array(27)(19),
      output(28) => mem_array(28)(19),
      output(29) => mem_array(29)(19),
      output(30) => mem_array(30)(19),
      output(31) => mem_array(31)(19),
      output(32) => mem_array(32)(19),
      output(33) => mem_array(33)(19),
      output(34) => mem_array(34)(19),
      output(35) => mem_array(35)(19)
      );
  rom20 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000010100000000010000011100000000")
    port map (
      enable_o   => mem_enable_lines(20),
      output(0)  => mem_array(0)(20),
      output(1)  => mem_array(1)(20),
      output(2)  => mem_array(2)(20),
      output(3)  => mem_array(3)(20),
      output(4)  => mem_array(4)(20),
      output(5)  => mem_array(5)(20),
      output(6)  => mem_array(6)(20),
      output(7)  => mem_array(7)(20),
      output(8)  => mem_array(8)(20),
      output(9)  => mem_array(9)(20),
      output(10) => mem_array(10)(20),
      output(11) => mem_array(11)(20),
      output(12) => mem_array(12)(20),
      output(13) => mem_array(13)(20),
      output(14) => mem_array(14)(20),
      output(15) => mem_array(15)(20),
      output(16) => mem_array(16)(20),
      output(17) => mem_array(17)(20),
      output(18) => mem_array(18)(20),
      output(19) => mem_array(19)(20),
      output(20) => mem_array(20)(20),
      output(21) => mem_array(21)(20),
      output(22) => mem_array(22)(20),
      output(23) => mem_array(23)(20),
      output(24) => mem_array(24)(20),
      output(25) => mem_array(25)(20),
      output(26) => mem_array(26)(20),
      output(27) => mem_array(27)(20),
      output(28) => mem_array(28)(20),
      output(29) => mem_array(29)(20),
      output(30) => mem_array(30)(20),
      output(31) => mem_array(31)(20),
      output(32) => mem_array(32)(20),
      output(33) => mem_array(33)(20),
      output(34) => mem_array(34)(20),
      output(35) => mem_array(35)(20)
      );
  rom21 : entity work.rom
    generic map (
      bits  => 36,
      value => "101000000011011000000000110001000000")
    port map (
      enable_o   => mem_enable_lines(21),
      output(0)  => mem_array(0)(21),
      output(1)  => mem_array(1)(21),
      output(2)  => mem_array(2)(21),
      output(3)  => mem_array(3)(21),
      output(4)  => mem_array(4)(21),
      output(5)  => mem_array(5)(21),
      output(6)  => mem_array(6)(21),
      output(7)  => mem_array(7)(21),
      output(8)  => mem_array(8)(21),
      output(9)  => mem_array(9)(21),
      output(10) => mem_array(10)(21),
      output(11) => mem_array(11)(21),
      output(12) => mem_array(12)(21),
      output(13) => mem_array(13)(21),
      output(14) => mem_array(14)(21),
      output(15) => mem_array(15)(21),
      output(16) => mem_array(16)(21),
      output(17) => mem_array(17)(21),
      output(18) => mem_array(18)(21),
      output(19) => mem_array(19)(21),
      output(20) => mem_array(20)(21),
      output(21) => mem_array(21)(21),
      output(22) => mem_array(22)(21),
      output(23) => mem_array(23)(21),
      output(24) => mem_array(24)(21),
      output(25) => mem_array(25)(21),
      output(26) => mem_array(26)(21),
      output(27) => mem_array(27)(21),
      output(28) => mem_array(28)(21),
      output(29) => mem_array(29)(21),
      output(30) => mem_array(30)(21),
      output(31) => mem_array(31)(21),
      output(32) => mem_array(32)(21),
      output(33) => mem_array(33)(21),
      output(34) => mem_array(34)(21),
      output(35) => mem_array(35)(21)
      );
  rom22 : entity work.rom
    generic map (
      bits  => 36,
      value => "000100111000001101010000001000010001")
    port map (
      enable_o   => mem_enable_lines(22),
      output(0)  => mem_array(0)(22),
      output(1)  => mem_array(1)(22),
      output(2)  => mem_array(2)(22),
      output(3)  => mem_array(3)(22),
      output(4)  => mem_array(4)(22),
      output(5)  => mem_array(5)(22),
      output(6)  => mem_array(6)(22),
      output(7)  => mem_array(7)(22),
      output(8)  => mem_array(8)(22),
      output(9)  => mem_array(9)(22),
      output(10) => mem_array(10)(22),
      output(11) => mem_array(11)(22),
      output(12) => mem_array(12)(22),
      output(13) => mem_array(13)(22),
      output(14) => mem_array(14)(22),
      output(15) => mem_array(15)(22),
      output(16) => mem_array(16)(22),
      output(17) => mem_array(17)(22),
      output(18) => mem_array(18)(22),
      output(19) => mem_array(19)(22),
      output(20) => mem_array(20)(22),
      output(21) => mem_array(21)(22),
      output(22) => mem_array(22)(22),
      output(23) => mem_array(23)(22),
      output(24) => mem_array(24)(22),
      output(25) => mem_array(25)(22),
      output(26) => mem_array(26)(22),
      output(27) => mem_array(27)(22),
      output(28) => mem_array(28)(22),
      output(29) => mem_array(29)(22),
      output(30) => mem_array(30)(22),
      output(31) => mem_array(31)(22),
      output(32) => mem_array(32)(22),
      output(33) => mem_array(33)(22),
      output(34) => mem_array(34)(22),
      output(35) => mem_array(35)(22)
      );
  rom23 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000001000000011000001000000000")
    port map (
      enable_o   => mem_enable_lines(23),
      output(0)  => mem_array(0)(23),
      output(1)  => mem_array(1)(23),
      output(2)  => mem_array(2)(23),
      output(3)  => mem_array(3)(23),
      output(4)  => mem_array(4)(23),
      output(5)  => mem_array(5)(23),
      output(6)  => mem_array(6)(23),
      output(7)  => mem_array(7)(23),
      output(8)  => mem_array(8)(23),
      output(9)  => mem_array(9)(23),
      output(10) => mem_array(10)(23),
      output(11) => mem_array(11)(23),
      output(12) => mem_array(12)(23),
      output(13) => mem_array(13)(23),
      output(14) => mem_array(14)(23),
      output(15) => mem_array(15)(23),
      output(16) => mem_array(16)(23),
      output(17) => mem_array(17)(23),
      output(18) => mem_array(18)(23),
      output(19) => mem_array(19)(23),
      output(20) => mem_array(20)(23),
      output(21) => mem_array(21)(23),
      output(22) => mem_array(22)(23),
      output(23) => mem_array(23)(23),
      output(24) => mem_array(24)(23),
      output(25) => mem_array(25)(23),
      output(26) => mem_array(26)(23),
      output(27) => mem_array(27)(23),
      output(28) => mem_array(28)(23),
      output(29) => mem_array(29)(23),
      output(30) => mem_array(30)(23),
      output(31) => mem_array(31)(23),
      output(32) => mem_array(32)(23),
      output(33) => mem_array(33)(23),
      output(34) => mem_array(34)(23),
      output(35) => mem_array(35)(23)
      );
  rom24 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000110000000001010010000000")
    port map (
      enable_o   => mem_enable_lines(24),
      output(0)  => mem_array(0)(24),
      output(1)  => mem_array(1)(24),
      output(2)  => mem_array(2)(24),
      output(3)  => mem_array(3)(24),
      output(4)  => mem_array(4)(24),
      output(5)  => mem_array(5)(24),
      output(6)  => mem_array(6)(24),
      output(7)  => mem_array(7)(24),
      output(8)  => mem_array(8)(24),
      output(9)  => mem_array(9)(24),
      output(10) => mem_array(10)(24),
      output(11) => mem_array(11)(24),
      output(12) => mem_array(12)(24),
      output(13) => mem_array(13)(24),
      output(14) => mem_array(14)(24),
      output(15) => mem_array(15)(24),
      output(16) => mem_array(16)(24),
      output(17) => mem_array(17)(24),
      output(18) => mem_array(18)(24),
      output(19) => mem_array(19)(24),
      output(20) => mem_array(20)(24),
      output(21) => mem_array(21)(24),
      output(22) => mem_array(22)(24),
      output(23) => mem_array(23)(24),
      output(24) => mem_array(24)(24),
      output(25) => mem_array(25)(24),
      output(26) => mem_array(26)(24),
      output(27) => mem_array(27)(24),
      output(28) => mem_array(28)(24),
      output(29) => mem_array(29)(24),
      output(30) => mem_array(30)(24),
      output(31) => mem_array(31)(24),
      output(32) => mem_array(32)(24),
      output(33) => mem_array(33)(24),
      output(34) => mem_array(34)(24),
      output(35) => mem_array(35)(24)
      );
  rom25 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001010000000010111000001101010000")
    port map (
      enable_o   => mem_enable_lines(25),
      output(0)  => mem_array(0)(25),
      output(1)  => mem_array(1)(25),
      output(2)  => mem_array(2)(25),
      output(3)  => mem_array(3)(25),
      output(4)  => mem_array(4)(25),
      output(5)  => mem_array(5)(25),
      output(6)  => mem_array(6)(25),
      output(7)  => mem_array(7)(25),
      output(8)  => mem_array(8)(25),
      output(9)  => mem_array(9)(25),
      output(10) => mem_array(10)(25),
      output(11) => mem_array(11)(25),
      output(12) => mem_array(12)(25),
      output(13) => mem_array(13)(25),
      output(14) => mem_array(14)(25),
      output(15) => mem_array(15)(25),
      output(16) => mem_array(16)(25),
      output(17) => mem_array(17)(25),
      output(18) => mem_array(18)(25),
      output(19) => mem_array(19)(25),
      output(20) => mem_array(20)(25),
      output(21) => mem_array(21)(25),
      output(22) => mem_array(22)(25),
      output(23) => mem_array(23)(25),
      output(24) => mem_array(24)(25),
      output(25) => mem_array(25)(25),
      output(26) => mem_array(26)(25),
      output(27) => mem_array(27)(25),
      output(28) => mem_array(28)(25),
      output(29) => mem_array(29)(25),
      output(30) => mem_array(30)(25),
      output(31) => mem_array(31)(25),
      output(32) => mem_array(32)(25),
      output(33) => mem_array(33)(25),
      output(34) => mem_array(34)(25),
      output(35) => mem_array(35)(25)
      );
  rom26 : entity work.rom
    generic map (
      bits  => 36,
      value => "001000010001000000000001000000010100")
    port map (
      enable_o   => mem_enable_lines(26),
      output(0)  => mem_array(0)(26),
      output(1)  => mem_array(1)(26),
      output(2)  => mem_array(2)(26),
      output(3)  => mem_array(3)(26),
      output(4)  => mem_array(4)(26),
      output(5)  => mem_array(5)(26),
      output(6)  => mem_array(6)(26),
      output(7)  => mem_array(7)(26),
      output(8)  => mem_array(8)(26),
      output(9)  => mem_array(9)(26),
      output(10) => mem_array(10)(26),
      output(11) => mem_array(11)(26),
      output(12) => mem_array(12)(26),
      output(13) => mem_array(13)(26),
      output(14) => mem_array(14)(26),
      output(15) => mem_array(15)(26),
      output(16) => mem_array(16)(26),
      output(17) => mem_array(17)(26),
      output(18) => mem_array(18)(26),
      output(19) => mem_array(19)(26),
      output(20) => mem_array(20)(26),
      output(21) => mem_array(21)(26),
      output(22) => mem_array(22)(26),
      output(23) => mem_array(23)(26),
      output(24) => mem_array(24)(26),
      output(25) => mem_array(25)(26),
      output(26) => mem_array(26)(26),
      output(27) => mem_array(27)(26),
      output(28) => mem_array(28)(26),
      output(29) => mem_array(29)(26),
      output(30) => mem_array(30)(26),
      output(31) => mem_array(31)(26),
      output(32) => mem_array(32)(26),
      output(33) => mem_array(33)(26),
      output(34) => mem_array(34)(26),
      output(35) => mem_array(35)(26)
      );
  rom27 : entity work.rom
    generic map (
      bits  => 36,
      value => "001000010100001000000000110010000011")
    port map (
      enable_o   => mem_enable_lines(27),
      output(0)  => mem_array(0)(27),
      output(1)  => mem_array(1)(27),
      output(2)  => mem_array(2)(27),
      output(3)  => mem_array(3)(27),
      output(4)  => mem_array(4)(27),
      output(5)  => mem_array(5)(27),
      output(6)  => mem_array(6)(27),
      output(7)  => mem_array(7)(27),
      output(8)  => mem_array(8)(27),
      output(9)  => mem_array(9)(27),
      output(10) => mem_array(10)(27),
      output(11) => mem_array(11)(27),
      output(12) => mem_array(12)(27),
      output(13) => mem_array(13)(27),
      output(14) => mem_array(14)(27),
      output(15) => mem_array(15)(27),
      output(16) => mem_array(16)(27),
      output(17) => mem_array(17)(27),
      output(18) => mem_array(18)(27),
      output(19) => mem_array(19)(27),
      output(20) => mem_array(20)(27),
      output(21) => mem_array(21)(27),
      output(22) => mem_array(22)(27),
      output(23) => mem_array(23)(27),
      output(24) => mem_array(24)(27),
      output(25) => mem_array(25)(27),
      output(26) => mem_array(26)(27),
      output(27) => mem_array(27)(27),
      output(28) => mem_array(28)(27),
      output(29) => mem_array(29)(27),
      output(30) => mem_array(30)(27),
      output(31) => mem_array(31)(27),
      output(32) => mem_array(32)(27),
      output(33) => mem_array(33)(27),
      output(34) => mem_array(34)(27),
      output(35) => mem_array(35)(27)
      );
  rom28 : entity work.rom
    generic map (
      bits  => 36,
      value => "110000000000101000110000000011010000")
    port map (
      enable_o   => mem_enable_lines(28),
      output(0)  => mem_array(0)(28),
      output(1)  => mem_array(1)(28),
      output(2)  => mem_array(2)(28),
      output(3)  => mem_array(3)(28),
      output(4)  => mem_array(4)(28),
      output(5)  => mem_array(5)(28),
      output(6)  => mem_array(6)(28),
      output(7)  => mem_array(7)(28),
      output(8)  => mem_array(8)(28),
      output(9)  => mem_array(9)(28),
      output(10) => mem_array(10)(28),
      output(11) => mem_array(11)(28),
      output(12) => mem_array(12)(28),
      output(13) => mem_array(13)(28),
      output(14) => mem_array(14)(28),
      output(15) => mem_array(15)(28),
      output(16) => mem_array(16)(28),
      output(17) => mem_array(17)(28),
      output(18) => mem_array(18)(28),
      output(19) => mem_array(19)(28),
      output(20) => mem_array(20)(28),
      output(21) => mem_array(21)(28),
      output(22) => mem_array(22)(28),
      output(23) => mem_array(23)(28),
      output(24) => mem_array(24)(28),
      output(25) => mem_array(25)(28),
      output(26) => mem_array(26)(28),
      output(27) => mem_array(27)(28),
      output(28) => mem_array(28)(28),
      output(29) => mem_array(29)(28),
      output(30) => mem_array(30)(28),
      output(31) => mem_array(31)(28),
      output(32) => mem_array(32)(28),
      output(33) => mem_array(33)(28),
      output(34) => mem_array(34)(28),
      output(35) => mem_array(35)(28)
      );
  rom29 : entity work.rom
    generic map (
      bits  => 36,
      value => "001101010000010010000100000000001101")
    port map (
      enable_o   => mem_enable_lines(29),
      output(0)  => mem_array(0)(29),
      output(1)  => mem_array(1)(29),
      output(2)  => mem_array(2)(29),
      output(3)  => mem_array(3)(29),
      output(4)  => mem_array(4)(29),
      output(5)  => mem_array(5)(29),
      output(6)  => mem_array(6)(29),
      output(7)  => mem_array(7)(29),
      output(8)  => mem_array(8)(29),
      output(9)  => mem_array(9)(29),
      output(10) => mem_array(10)(29),
      output(11) => mem_array(11)(29),
      output(12) => mem_array(12)(29),
      output(13) => mem_array(13)(29),
      output(14) => mem_array(14)(29),
      output(15) => mem_array(15)(29),
      output(16) => mem_array(16)(29),
      output(17) => mem_array(17)(29),
      output(18) => mem_array(18)(29),
      output(19) => mem_array(19)(29),
      output(20) => mem_array(20)(29),
      output(21) => mem_array(21)(29),
      output(22) => mem_array(22)(29),
      output(23) => mem_array(23)(29),
      output(24) => mem_array(24)(29),
      output(25) => mem_array(25)(29),
      output(26) => mem_array(26)(29),
      output(27) => mem_array(27)(29),
      output(28) => mem_array(28)(29),
      output(29) => mem_array(29)(29),
      output(30) => mem_array(30)(29),
      output(31) => mem_array(31)(29),
      output(32) => mem_array(32)(29),
      output(33) => mem_array(33)(29),
      output(34) => mem_array(34)(29),
      output(35) => mem_array(35)(29)
      );
  rom30 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000110101000000100101000100000000")
    port map (
      enable_o   => mem_enable_lines(30),
      output(0)  => mem_array(0)(30),
      output(1)  => mem_array(1)(30),
      output(2)  => mem_array(2)(30),
      output(3)  => mem_array(3)(30),
      output(4)  => mem_array(4)(30),
      output(5)  => mem_array(5)(30),
      output(6)  => mem_array(6)(30),
      output(7)  => mem_array(7)(30),
      output(8)  => mem_array(8)(30),
      output(9)  => mem_array(9)(30),
      output(10) => mem_array(10)(30),
      output(11) => mem_array(11)(30),
      output(12) => mem_array(12)(30),
      output(13) => mem_array(13)(30),
      output(14) => mem_array(14)(30),
      output(15) => mem_array(15)(30),
      output(16) => mem_array(16)(30),
      output(17) => mem_array(17)(30),
      output(18) => mem_array(18)(30),
      output(19) => mem_array(19)(30),
      output(20) => mem_array(20)(30),
      output(21) => mem_array(21)(30),
      output(22) => mem_array(22)(30),
      output(23) => mem_array(23)(30),
      output(24) => mem_array(24)(30),
      output(25) => mem_array(25)(30),
      output(26) => mem_array(26)(30),
      output(27) => mem_array(27)(30),
      output(28) => mem_array(28)(30),
      output(29) => mem_array(29)(30),
      output(30) => mem_array(30)(30),
      output(31) => mem_array(31)(30),
      output(32) => mem_array(32)(30),
      output(33) => mem_array(33)(30),
      output(34) => mem_array(34)(30),
      output(35) => mem_array(35)(30)
      );
  rom31 : entity work.rom
    generic map (
      bits  => 36,
      value => "000100000001010000100000000000000000")
    port map (
      enable_o   => mem_enable_lines(31),
      output(0)  => mem_array(0)(31),
      output(1)  => mem_array(1)(31),
      output(2)  => mem_array(2)(31),
      output(3)  => mem_array(3)(31),
      output(4)  => mem_array(4)(31),
      output(5)  => mem_array(5)(31),
      output(6)  => mem_array(6)(31),
      output(7)  => mem_array(7)(31),
      output(8)  => mem_array(8)(31),
      output(9)  => mem_array(9)(31),
      output(10) => mem_array(10)(31),
      output(11) => mem_array(11)(31),
      output(12) => mem_array(12)(31),
      output(13) => mem_array(13)(31),
      output(14) => mem_array(14)(31),
      output(15) => mem_array(15)(31),
      output(16) => mem_array(16)(31),
      output(17) => mem_array(17)(31),
      output(18) => mem_array(18)(31),
      output(19) => mem_array(19)(31),
      output(20) => mem_array(20)(31),
      output(21) => mem_array(21)(31),
      output(22) => mem_array(22)(31),
      output(23) => mem_array(23)(31),
      output(24) => mem_array(24)(31),
      output(25) => mem_array(25)(31),
      output(26) => mem_array(26)(31),
      output(27) => mem_array(27)(31),
      output(28) => mem_array(28)(31),
      output(29) => mem_array(29)(31),
      output(30) => mem_array(30)(31),
      output(31) => mem_array(31)(31),
      output(32) => mem_array(32)(31),
      output(33) => mem_array(33)(31),
      output(34) => mem_array(34)(31),
      output(35) => mem_array(35)(31)
      );
  rom32 : entity work.rom
    generic map (
      bits  => 36,
      value => "000011101000001111000000000010000011")
    port map (
      enable_o   => mem_enable_lines(32),
      output(0)  => mem_array(0)(32),
      output(1)  => mem_array(1)(32),
      output(2)  => mem_array(2)(32),
      output(3)  => mem_array(3)(32),
      output(4)  => mem_array(4)(32),
      output(5)  => mem_array(5)(32),
      output(6)  => mem_array(6)(32),
      output(7)  => mem_array(7)(32),
      output(8)  => mem_array(8)(32),
      output(9)  => mem_array(9)(32),
      output(10) => mem_array(10)(32),
      output(11) => mem_array(11)(32),
      output(12) => mem_array(12)(32),
      output(13) => mem_array(13)(32),
      output(14) => mem_array(14)(32),
      output(15) => mem_array(15)(32),
      output(16) => mem_array(16)(32),
      output(17) => mem_array(17)(32),
      output(18) => mem_array(18)(32),
      output(19) => mem_array(19)(32),
      output(20) => mem_array(20)(32),
      output(21) => mem_array(21)(32),
      output(22) => mem_array(22)(32),
      output(23) => mem_array(23)(32),
      output(24) => mem_array(24)(32),
      output(25) => mem_array(25)(32),
      output(26) => mem_array(26)(32),
      output(27) => mem_array(27)(32),
      output(28) => mem_array(28)(32),
      output(29) => mem_array(29)(32),
      output(30) => mem_array(30)(32),
      output(31) => mem_array(31)(32),
      output(32) => mem_array(32)(32),
      output(33) => mem_array(33)(32),
      output(34) => mem_array(34)(32),
      output(35) => mem_array(35)(32)
      );
  rom33 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001111000000010100000000010100")
    port map (
      enable_o   => mem_enable_lines(33),
      output(0)  => mem_array(0)(33),
      output(1)  => mem_array(1)(33),
      output(2)  => mem_array(2)(33),
      output(3)  => mem_array(3)(33),
      output(4)  => mem_array(4)(33),
      output(5)  => mem_array(5)(33),
      output(6)  => mem_array(6)(33),
      output(7)  => mem_array(7)(33),
      output(8)  => mem_array(8)(33),
      output(9)  => mem_array(9)(33),
      output(10) => mem_array(10)(33),
      output(11) => mem_array(11)(33),
      output(12) => mem_array(12)(33),
      output(13) => mem_array(13)(33),
      output(14) => mem_array(14)(33),
      output(15) => mem_array(15)(33),
      output(16) => mem_array(16)(33),
      output(17) => mem_array(17)(33),
      output(18) => mem_array(18)(33),
      output(19) => mem_array(19)(33),
      output(20) => mem_array(20)(33),
      output(21) => mem_array(21)(33),
      output(22) => mem_array(22)(33),
      output(23) => mem_array(23)(33),
      output(24) => mem_array(24)(33),
      output(25) => mem_array(25)(33),
      output(26) => mem_array(26)(33),
      output(27) => mem_array(27)(33),
      output(28) => mem_array(28)(33),
      output(29) => mem_array(29)(33),
      output(30) => mem_array(30)(33),
      output(31) => mem_array(31)(33),
      output(32) => mem_array(32)(33),
      output(33) => mem_array(33)(33),
      output(34) => mem_array(34)(33),
      output(35) => mem_array(35)(33)
      );
  rom34 : entity work.rom
    generic map (
      bits  => 36,
      value => "011100000000111110000011011000000100")
    port map (
      enable_o   => mem_enable_lines(34),
      output(0)  => mem_array(0)(34),
      output(1)  => mem_array(1)(34),
      output(2)  => mem_array(2)(34),
      output(3)  => mem_array(3)(34),
      output(4)  => mem_array(4)(34),
      output(5)  => mem_array(5)(34),
      output(6)  => mem_array(6)(34),
      output(7)  => mem_array(7)(34),
      output(8)  => mem_array(8)(34),
      output(9)  => mem_array(9)(34),
      output(10) => mem_array(10)(34),
      output(11) => mem_array(11)(34),
      output(12) => mem_array(12)(34),
      output(13) => mem_array(13)(34),
      output(14) => mem_array(14)(34),
      output(15) => mem_array(15)(34),
      output(16) => mem_array(16)(34),
      output(17) => mem_array(17)(34),
      output(18) => mem_array(18)(34),
      output(19) => mem_array(19)(34),
      output(20) => mem_array(20)(34),
      output(21) => mem_array(21)(34),
      output(22) => mem_array(22)(34),
      output(23) => mem_array(23)(34),
      output(24) => mem_array(24)(34),
      output(25) => mem_array(25)(34),
      output(26) => mem_array(26)(34),
      output(27) => mem_array(27)(34),
      output(28) => mem_array(28)(34),
      output(29) => mem_array(29)(34),
      output(30) => mem_array(30)(34),
      output(31) => mem_array(31)(34),
      output(32) => mem_array(32)(34),
      output(33) => mem_array(33)(34),
      output(34) => mem_array(34)(34),
      output(35) => mem_array(35)(34)
      );
  rom35 : entity work.rom
    generic map (
      bits  => 36,
      value => "101001000000000100000000001101010000")
    port map (
      enable_o   => mem_enable_lines(35),
      output(0)  => mem_array(0)(35),
      output(1)  => mem_array(1)(35),
      output(2)  => mem_array(2)(35),
      output(3)  => mem_array(3)(35),
      output(4)  => mem_array(4)(35),
      output(5)  => mem_array(5)(35),
      output(6)  => mem_array(6)(35),
      output(7)  => mem_array(7)(35),
      output(8)  => mem_array(8)(35),
      output(9)  => mem_array(9)(35),
      output(10) => mem_array(10)(35),
      output(11) => mem_array(11)(35),
      output(12) => mem_array(12)(35),
      output(13) => mem_array(13)(35),
      output(14) => mem_array(14)(35),
      output(15) => mem_array(15)(35),
      output(16) => mem_array(16)(35),
      output(17) => mem_array(17)(35),
      output(18) => mem_array(18)(35),
      output(19) => mem_array(19)(35),
      output(20) => mem_array(20)(35),
      output(21) => mem_array(21)(35),
      output(22) => mem_array(22)(35),
      output(23) => mem_array(23)(35),
      output(24) => mem_array(24)(35),
      output(25) => mem_array(25)(35),
      output(26) => mem_array(26)(35),
      output(27) => mem_array(27)(35),
      output(28) => mem_array(28)(35),
      output(29) => mem_array(29)(35),
      output(30) => mem_array(30)(35),
      output(31) => mem_array(31)(35),
      output(32) => mem_array(32)(35),
      output(33) => mem_array(33)(35),
      output(34) => mem_array(34)(35),
      output(35) => mem_array(35)(35)
      );
  rom36 : entity work.rom
    generic map (
      bits  => 36,
      value => "001000010001000000000001000000010100")
    port map (
      enable_o   => mem_enable_lines(36),
      output(0)  => mem_array(0)(36),
      output(1)  => mem_array(1)(36),
      output(2)  => mem_array(2)(36),
      output(3)  => mem_array(3)(36),
      output(4)  => mem_array(4)(36),
      output(5)  => mem_array(5)(36),
      output(6)  => mem_array(6)(36),
      output(7)  => mem_array(7)(36),
      output(8)  => mem_array(8)(36),
      output(9)  => mem_array(9)(36),
      output(10) => mem_array(10)(36),
      output(11) => mem_array(11)(36),
      output(12) => mem_array(12)(36),
      output(13) => mem_array(13)(36),
      output(14) => mem_array(14)(36),
      output(15) => mem_array(15)(36),
      output(16) => mem_array(16)(36),
      output(17) => mem_array(17)(36),
      output(18) => mem_array(18)(36),
      output(19) => mem_array(19)(36),
      output(20) => mem_array(20)(36),
      output(21) => mem_array(21)(36),
      output(22) => mem_array(22)(36),
      output(23) => mem_array(23)(36),
      output(24) => mem_array(24)(36),
      output(25) => mem_array(25)(36),
      output(26) => mem_array(26)(36),
      output(27) => mem_array(27)(36),
      output(28) => mem_array(28)(36),
      output(29) => mem_array(29)(36),
      output(30) => mem_array(30)(36),
      output(31) => mem_array(31)(36),
      output(32) => mem_array(32)(36),
      output(33) => mem_array(33)(36),
      output(34) => mem_array(34)(36),
      output(35) => mem_array(35)(36)
      );
  rom37 : entity work.rom
    generic map (
      bits  => 36,
      value => "001000000000000000000001000100001001")
    port map (
      enable_o   => mem_enable_lines(37),
      output(0)  => mem_array(0)(37),
      output(1)  => mem_array(1)(37),
      output(2)  => mem_array(2)(37),
      output(3)  => mem_array(3)(37),
      output(4)  => mem_array(4)(37),
      output(5)  => mem_array(5)(37),
      output(6)  => mem_array(6)(37),
      output(7)  => mem_array(7)(37),
      output(8)  => mem_array(8)(37),
      output(9)  => mem_array(9)(37),
      output(10) => mem_array(10)(37),
      output(11) => mem_array(11)(37),
      output(12) => mem_array(12)(37),
      output(13) => mem_array(13)(37),
      output(14) => mem_array(14)(37),
      output(15) => mem_array(15)(37),
      output(16) => mem_array(16)(37),
      output(17) => mem_array(17)(37),
      output(18) => mem_array(18)(37),
      output(19) => mem_array(19)(37),
      output(20) => mem_array(20)(37),
      output(21) => mem_array(21)(37),
      output(22) => mem_array(22)(37),
      output(23) => mem_array(23)(37),
      output(24) => mem_array(24)(37),
      output(25) => mem_array(25)(37),
      output(26) => mem_array(26)(37),
      output(27) => mem_array(27)(37),
      output(28) => mem_array(28)(37),
      output(29) => mem_array(29)(37),
      output(30) => mem_array(30)(37),
      output(31) => mem_array(31)(37),
      output(32) => mem_array(32)(37),
      output(33) => mem_array(33)(37),
      output(34) => mem_array(34)(37),
      output(35) => mem_array(35)(37)
      );
  rom38 : entity work.rom
    generic map (
      bits  => 36,
      value => "010010000000000000110000000100011000")
    port map (
      enable_o   => mem_enable_lines(38),
      output(0)  => mem_array(0)(38),
      output(1)  => mem_array(1)(38),
      output(2)  => mem_array(2)(38),
      output(3)  => mem_array(3)(38),
      output(4)  => mem_array(4)(38),
      output(5)  => mem_array(5)(38),
      output(6)  => mem_array(6)(38),
      output(7)  => mem_array(7)(38),
      output(8)  => mem_array(8)(38),
      output(9)  => mem_array(9)(38),
      output(10) => mem_array(10)(38),
      output(11) => mem_array(11)(38),
      output(12) => mem_array(12)(38),
      output(13) => mem_array(13)(38),
      output(14) => mem_array(14)(38),
      output(15) => mem_array(15)(38),
      output(16) => mem_array(16)(38),
      output(17) => mem_array(17)(38),
      output(18) => mem_array(18)(38),
      output(19) => mem_array(19)(38),
      output(20) => mem_array(20)(38),
      output(21) => mem_array(21)(38),
      output(22) => mem_array(22)(38),
      output(23) => mem_array(23)(38),
      output(24) => mem_array(24)(38),
      output(25) => mem_array(25)(38),
      output(26) => mem_array(26)(38),
      output(27) => mem_array(27)(38),
      output(28) => mem_array(28)(38),
      output(29) => mem_array(29)(38),
      output(30) => mem_array(30)(38),
      output(31) => mem_array(31)(38),
      output(32) => mem_array(32)(38),
      output(33) => mem_array(33)(38),
      output(34) => mem_array(34)(38),
      output(35) => mem_array(35)(38)
      );
  rom39 : entity work.rom
    generic map (
      bits  => 36,
      value => "000111001000000000000011000000001100")
    port map (
      enable_o   => mem_enable_lines(39),
      output(0)  => mem_array(0)(39),
      output(1)  => mem_array(1)(39),
      output(2)  => mem_array(2)(39),
      output(3)  => mem_array(3)(39),
      output(4)  => mem_array(4)(39),
      output(5)  => mem_array(5)(39),
      output(6)  => mem_array(6)(39),
      output(7)  => mem_array(7)(39),
      output(8)  => mem_array(8)(39),
      output(9)  => mem_array(9)(39),
      output(10) => mem_array(10)(39),
      output(11) => mem_array(11)(39),
      output(12) => mem_array(12)(39),
      output(13) => mem_array(13)(39),
      output(14) => mem_array(14)(39),
      output(15) => mem_array(15)(39),
      output(16) => mem_array(16)(39),
      output(17) => mem_array(17)(39),
      output(18) => mem_array(18)(39),
      output(19) => mem_array(19)(39),
      output(20) => mem_array(20)(39),
      output(21) => mem_array(21)(39),
      output(22) => mem_array(22)(39),
      output(23) => mem_array(23)(39),
      output(24) => mem_array(24)(39),
      output(25) => mem_array(25)(39),
      output(26) => mem_array(26)(39),
      output(27) => mem_array(27)(39),
      output(28) => mem_array(28)(39),
      output(29) => mem_array(29)(39),
      output(30) => mem_array(30)(39),
      output(31) => mem_array(31)(39),
      output(32) => mem_array(32)(39),
      output(33) => mem_array(33)(39),
      output(34) => mem_array(34)(39),
      output(35) => mem_array(35)(39)
      );
  rom40 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000111100000000001010010100000001")
    port map (
      enable_o   => mem_enable_lines(40),
      output(0)  => mem_array(0)(40),
      output(1)  => mem_array(1)(40),
      output(2)  => mem_array(2)(40),
      output(3)  => mem_array(3)(40),
      output(4)  => mem_array(4)(40),
      output(5)  => mem_array(5)(40),
      output(6)  => mem_array(6)(40),
      output(7)  => mem_array(7)(40),
      output(8)  => mem_array(8)(40),
      output(9)  => mem_array(9)(40),
      output(10) => mem_array(10)(40),
      output(11) => mem_array(11)(40),
      output(12) => mem_array(12)(40),
      output(13) => mem_array(13)(40),
      output(14) => mem_array(14)(40),
      output(15) => mem_array(15)(40),
      output(16) => mem_array(16)(40),
      output(17) => mem_array(17)(40),
      output(18) => mem_array(18)(40),
      output(19) => mem_array(19)(40),
      output(20) => mem_array(20)(40),
      output(21) => mem_array(21)(40),
      output(22) => mem_array(22)(40),
      output(23) => mem_array(23)(40),
      output(24) => mem_array(24)(40),
      output(25) => mem_array(25)(40),
      output(26) => mem_array(26)(40),
      output(27) => mem_array(27)(40),
      output(28) => mem_array(28)(40),
      output(29) => mem_array(29)(40),
      output(30) => mem_array(30)(40),
      output(31) => mem_array(31)(40),
      output(32) => mem_array(32)(40),
      output(33) => mem_array(33)(40),
      output(34) => mem_array(34)(40),
      output(35) => mem_array(35)(40)
      );
  rom41 : entity work.rom
    generic map (
      bits  => 36,
      value => "001010001001010010000000000000110000")
    port map (
      enable_o   => mem_enable_lines(41),
      output(0)  => mem_array(0)(41),
      output(1)  => mem_array(1)(41),
      output(2)  => mem_array(2)(41),
      output(3)  => mem_array(3)(41),
      output(4)  => mem_array(4)(41),
      output(5)  => mem_array(5)(41),
      output(6)  => mem_array(6)(41),
      output(7)  => mem_array(7)(41),
      output(8)  => mem_array(8)(41),
      output(9)  => mem_array(9)(41),
      output(10) => mem_array(10)(41),
      output(11) => mem_array(11)(41),
      output(12) => mem_array(12)(41),
      output(13) => mem_array(13)(41),
      output(14) => mem_array(14)(41),
      output(15) => mem_array(15)(41),
      output(16) => mem_array(16)(41),
      output(17) => mem_array(17)(41),
      output(18) => mem_array(18)(41),
      output(19) => mem_array(19)(41),
      output(20) => mem_array(20)(41),
      output(21) => mem_array(21)(41),
      output(22) => mem_array(22)(41),
      output(23) => mem_array(23)(41),
      output(24) => mem_array(24)(41),
      output(25) => mem_array(25)(41),
      output(26) => mem_array(26)(41),
      output(27) => mem_array(27)(41),
      output(28) => mem_array(28)(41),
      output(29) => mem_array(29)(41),
      output(30) => mem_array(30)(41),
      output(31) => mem_array(31)(41),
      output(32) => mem_array(32)(41),
      output(33) => mem_array(33)(41),
      output(34) => mem_array(34)(41),
      output(35) => mem_array(35)(41)
      );
  rom42 : entity work.rom
    generic map (
      bits  => 36,
      value => "000100110000000111001000000000000011")
    port map (
      enable_o   => mem_enable_lines(42),
      output(0)  => mem_array(0)(42),
      output(1)  => mem_array(1)(42),
      output(2)  => mem_array(2)(42),
      output(3)  => mem_array(3)(42),
      output(4)  => mem_array(4)(42),
      output(5)  => mem_array(5)(42),
      output(6)  => mem_array(6)(42),
      output(7)  => mem_array(7)(42),
      output(8)  => mem_array(8)(42),
      output(9)  => mem_array(9)(42),
      output(10) => mem_array(10)(42),
      output(11) => mem_array(11)(42),
      output(12) => mem_array(12)(42),
      output(13) => mem_array(13)(42),
      output(14) => mem_array(14)(42),
      output(15) => mem_array(15)(42),
      output(16) => mem_array(16)(42),
      output(17) => mem_array(17)(42),
      output(18) => mem_array(18)(42),
      output(19) => mem_array(19)(42),
      output(20) => mem_array(20)(42),
      output(21) => mem_array(21)(42),
      output(22) => mem_array(22)(42),
      output(23) => mem_array(23)(42),
      output(24) => mem_array(24)(42),
      output(25) => mem_array(25)(42),
      output(26) => mem_array(26)(42),
      output(27) => mem_array(27)(42),
      output(28) => mem_array(28)(42),
      output(29) => mem_array(29)(42),
      output(30) => mem_array(30)(42),
      output(31) => mem_array(31)(42),
      output(32) => mem_array(32)(42),
      output(33) => mem_array(33)(42),
      output(34) => mem_array(34)(42),
      output(35) => mem_array(35)(42)
      );
  rom43 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001110100000111100000000001000")
    port map (
      enable_o   => mem_enable_lines(43),
      output(0)  => mem_array(0)(43),
      output(1)  => mem_array(1)(43),
      output(2)  => mem_array(2)(43),
      output(3)  => mem_array(3)(43),
      output(4)  => mem_array(4)(43),
      output(5)  => mem_array(5)(43),
      output(6)  => mem_array(6)(43),
      output(7)  => mem_array(7)(43),
      output(8)  => mem_array(8)(43),
      output(9)  => mem_array(9)(43),
      output(10) => mem_array(10)(43),
      output(11) => mem_array(11)(43),
      output(12) => mem_array(12)(43),
      output(13) => mem_array(13)(43),
      output(14) => mem_array(14)(43),
      output(15) => mem_array(15)(43),
      output(16) => mem_array(16)(43),
      output(17) => mem_array(17)(43),
      output(18) => mem_array(18)(43),
      output(19) => mem_array(19)(43),
      output(20) => mem_array(20)(43),
      output(21) => mem_array(21)(43),
      output(22) => mem_array(22)(43),
      output(23) => mem_array(23)(43),
      output(24) => mem_array(24)(43),
      output(25) => mem_array(25)(43),
      output(26) => mem_array(26)(43),
      output(27) => mem_array(27)(43),
      output(28) => mem_array(28)(43),
      output(29) => mem_array(29)(43),
      output(30) => mem_array(30)(43),
      output(31) => mem_array(31)(43),
      output(32) => mem_array(32)(43),
      output(33) => mem_array(33)(43),
      output(34) => mem_array(34)(43),
      output(35) => mem_array(35)(43)
      );
  rom44 : entity work.rom
    generic map (
      bits  => 36,
      value => "010100000001010000001001010010000000")
    port map (
      enable_o   => mem_enable_lines(44),
      output(0)  => mem_array(0)(44),
      output(1)  => mem_array(1)(44),
      output(2)  => mem_array(2)(44),
      output(3)  => mem_array(3)(44),
      output(4)  => mem_array(4)(44),
      output(5)  => mem_array(5)(44),
      output(6)  => mem_array(6)(44),
      output(7)  => mem_array(7)(44),
      output(8)  => mem_array(8)(44),
      output(9)  => mem_array(9)(44),
      output(10) => mem_array(10)(44),
      output(11) => mem_array(11)(44),
      output(12) => mem_array(12)(44),
      output(13) => mem_array(13)(44),
      output(14) => mem_array(14)(44),
      output(15) => mem_array(15)(44),
      output(16) => mem_array(16)(44),
      output(17) => mem_array(17)(44),
      output(18) => mem_array(18)(44),
      output(19) => mem_array(19)(44),
      output(20) => mem_array(20)(44),
      output(21) => mem_array(21)(44),
      output(22) => mem_array(22)(44),
      output(23) => mem_array(23)(44),
      output(24) => mem_array(24)(44),
      output(25) => mem_array(25)(44),
      output(26) => mem_array(26)(44),
      output(27) => mem_array(27)(44),
      output(28) => mem_array(28)(44),
      output(29) => mem_array(29)(44),
      output(30) => mem_array(30)(44),
      output(31) => mem_array(31)(44),
      output(32) => mem_array(32)(44),
      output(33) => mem_array(33)(44),
      output(34) => mem_array(34)(44),
      output(35) => mem_array(35)(44)
      );
  rom45 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000110000000101001000000111001000")
    port map (
      enable_o   => mem_enable_lines(45),
      output(0)  => mem_array(0)(45),
      output(1)  => mem_array(1)(45),
      output(2)  => mem_array(2)(45),
      output(3)  => mem_array(3)(45),
      output(4)  => mem_array(4)(45),
      output(5)  => mem_array(5)(45),
      output(6)  => mem_array(6)(45),
      output(7)  => mem_array(7)(45),
      output(8)  => mem_array(8)(45),
      output(9)  => mem_array(9)(45),
      output(10) => mem_array(10)(45),
      output(11) => mem_array(11)(45),
      output(12) => mem_array(12)(45),
      output(13) => mem_array(13)(45),
      output(14) => mem_array(14)(45),
      output(15) => mem_array(15)(45),
      output(16) => mem_array(16)(45),
      output(17) => mem_array(17)(45),
      output(18) => mem_array(18)(45),
      output(19) => mem_array(19)(45),
      output(20) => mem_array(20)(45),
      output(21) => mem_array(21)(45),
      output(22) => mem_array(22)(45),
      output(23) => mem_array(23)(45),
      output(24) => mem_array(24)(45),
      output(25) => mem_array(25)(45),
      output(26) => mem_array(26)(45),
      output(27) => mem_array(27)(45),
      output(28) => mem_array(28)(45),
      output(29) => mem_array(29)(45),
      output(30) => mem_array(30)(45),
      output(31) => mem_array(31)(45),
      output(32) => mem_array(32)(45),
      output(33) => mem_array(33)(45),
      output(34) => mem_array(34)(45),
      output(35) => mem_array(35)(45)
      );
  rom46 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000011000000001100100000111100")
    port map (
      enable_o   => mem_enable_lines(46),
      output(0)  => mem_array(0)(46),
      output(1)  => mem_array(1)(46),
      output(2)  => mem_array(2)(46),
      output(3)  => mem_array(3)(46),
      output(4)  => mem_array(4)(46),
      output(5)  => mem_array(5)(46),
      output(6)  => mem_array(6)(46),
      output(7)  => mem_array(7)(46),
      output(8)  => mem_array(8)(46),
      output(9)  => mem_array(9)(46),
      output(10) => mem_array(10)(46),
      output(11) => mem_array(11)(46),
      output(12) => mem_array(12)(46),
      output(13) => mem_array(13)(46),
      output(14) => mem_array(14)(46),
      output(15) => mem_array(15)(46),
      output(16) => mem_array(16)(46),
      output(17) => mem_array(17)(46),
      output(18) => mem_array(18)(46),
      output(19) => mem_array(19)(46),
      output(20) => mem_array(20)(46),
      output(21) => mem_array(21)(46),
      output(22) => mem_array(22)(46),
      output(23) => mem_array(23)(46),
      output(24) => mem_array(24)(46),
      output(25) => mem_array(25)(46),
      output(26) => mem_array(26)(46),
      output(27) => mem_array(27)(46),
      output(28) => mem_array(28)(46),
      output(29) => mem_array(29)(46),
      output(30) => mem_array(30)(46),
      output(31) => mem_array(31)(46),
      output(32) => mem_array(32)(46),
      output(33) => mem_array(33)(46),
      output(34) => mem_array(34)(46),
      output(35) => mem_array(35)(46)
      );
  rom47 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001010011000000001010110000011")
    port map (
      enable_o   => mem_enable_lines(47),
      output(0)  => mem_array(0)(47),
      output(1)  => mem_array(1)(47),
      output(2)  => mem_array(2)(47),
      output(3)  => mem_array(3)(47),
      output(4)  => mem_array(4)(47),
      output(5)  => mem_array(5)(47),
      output(6)  => mem_array(6)(47),
      output(7)  => mem_array(7)(47),
      output(8)  => mem_array(8)(47),
      output(9)  => mem_array(9)(47),
      output(10) => mem_array(10)(47),
      output(11) => mem_array(11)(47),
      output(12) => mem_array(12)(47),
      output(13) => mem_array(13)(47),
      output(14) => mem_array(14)(47),
      output(15) => mem_array(15)(47),
      output(16) => mem_array(16)(47),
      output(17) => mem_array(17)(47),
      output(18) => mem_array(18)(47),
      output(19) => mem_array(19)(47),
      output(20) => mem_array(20)(47),
      output(21) => mem_array(21)(47),
      output(22) => mem_array(22)(47),
      output(23) => mem_array(23)(47),
      output(24) => mem_array(24)(47),
      output(25) => mem_array(25)(47),
      output(26) => mem_array(26)(47),
      output(27) => mem_array(27)(47),
      output(28) => mem_array(28)(47),
      output(29) => mem_array(29)(47),
      output(30) => mem_array(30)(47),
      output(31) => mem_array(31)(47),
      output(32) => mem_array(32)(47),
      output(33) => mem_array(33)(47),
      output(34) => mem_array(34)(47),
      output(35) => mem_array(35)(47)
      );
  rom48 : entity work.rom
    generic map (
      bits  => 36,
      value => "110000000000101000110000000101100000")
    port map (
      enable_o   => mem_enable_lines(48),
      output(0)  => mem_array(0)(48),
      output(1)  => mem_array(1)(48),
      output(2)  => mem_array(2)(48),
      output(3)  => mem_array(3)(48),
      output(4)  => mem_array(4)(48),
      output(5)  => mem_array(5)(48),
      output(6)  => mem_array(6)(48),
      output(7)  => mem_array(7)(48),
      output(8)  => mem_array(8)(48),
      output(9)  => mem_array(9)(48),
      output(10) => mem_array(10)(48),
      output(11) => mem_array(11)(48),
      output(12) => mem_array(12)(48),
      output(13) => mem_array(13)(48),
      output(14) => mem_array(14)(48),
      output(15) => mem_array(15)(48),
      output(16) => mem_array(16)(48),
      output(17) => mem_array(17)(48),
      output(18) => mem_array(18)(48),
      output(19) => mem_array(19)(48),
      output(20) => mem_array(20)(48),
      output(21) => mem_array(21)(48),
      output(22) => mem_array(22)(48),
      output(23) => mem_array(23)(48),
      output(24) => mem_array(24)(48),
      output(25) => mem_array(25)(48),
      output(26) => mem_array(26)(48),
      output(27) => mem_array(27)(48),
      output(28) => mem_array(28)(48),
      output(29) => mem_array(29)(48),
      output(30) => mem_array(30)(48),
      output(31) => mem_array(31)(48),
      output(32) => mem_array(32)(48),
      output(33) => mem_array(33)(48),
      output(34) => mem_array(34)(48),
      output(35) => mem_array(35)(48)
      );
  rom49 : entity work.rom
    generic map (
      bits  => 36,
      value => "001101010000001000010001000000010110")
    port map (
      enable_o   => mem_enable_lines(49),
      output(0)  => mem_array(0)(49),
      output(1)  => mem_array(1)(49),
      output(2)  => mem_array(2)(49),
      output(3)  => mem_array(3)(49),
      output(4)  => mem_array(4)(49),
      output(5)  => mem_array(5)(49),
      output(6)  => mem_array(6)(49),
      output(7)  => mem_array(7)(49),
      output(8)  => mem_array(8)(49),
      output(9)  => mem_array(9)(49),
      output(10) => mem_array(10)(49),
      output(11) => mem_array(11)(49),
      output(12) => mem_array(12)(49),
      output(13) => mem_array(13)(49),
      output(14) => mem_array(14)(49),
      output(15) => mem_array(15)(49),
      output(16) => mem_array(16)(49),
      output(17) => mem_array(17)(49),
      output(18) => mem_array(18)(49),
      output(19) => mem_array(19)(49),
      output(20) => mem_array(20)(49),
      output(21) => mem_array(21)(49),
      output(22) => mem_array(22)(49),
      output(23) => mem_array(23)(49),
      output(24) => mem_array(24)(49),
      output(25) => mem_array(25)(49),
      output(26) => mem_array(26)(49),
      output(27) => mem_array(27)(49),
      output(28) => mem_array(28)(49),
      output(29) => mem_array(29)(49),
      output(30) => mem_array(30)(49),
      output(31) => mem_array(31)(49),
      output(32) => mem_array(32)(49),
      output(33) => mem_array(33)(49),
      output(34) => mem_array(34)(49),
      output(35) => mem_array(35)(49)
      );
  rom50 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000010100100000000000000000000001")
    port map (
      enable_o   => mem_enable_lines(50),
      output(0)  => mem_array(0)(50),
      output(1)  => mem_array(1)(50),
      output(2)  => mem_array(2)(50),
      output(3)  => mem_array(3)(50),
      output(4)  => mem_array(4)(50),
      output(5)  => mem_array(5)(50),
      output(6)  => mem_array(6)(50),
      output(7)  => mem_array(7)(50),
      output(8)  => mem_array(8)(50),
      output(9)  => mem_array(9)(50),
      output(10) => mem_array(10)(50),
      output(11) => mem_array(11)(50),
      output(12) => mem_array(12)(50),
      output(13) => mem_array(13)(50),
      output(14) => mem_array(14)(50),
      output(15) => mem_array(15)(50),
      output(16) => mem_array(16)(50),
      output(17) => mem_array(17)(50),
      output(18) => mem_array(18)(50),
      output(19) => mem_array(19)(50),
      output(20) => mem_array(20)(50),
      output(21) => mem_array(21)(50),
      output(22) => mem_array(22)(50),
      output(23) => mem_array(23)(50),
      output(24) => mem_array(24)(50),
      output(25) => mem_array(25)(50),
      output(26) => mem_array(26)(50),
      output(27) => mem_array(27)(50),
      output(28) => mem_array(28)(50),
      output(29) => mem_array(29)(50),
      output(30) => mem_array(30)(50),
      output(31) => mem_array(31)(50),
      output(32) => mem_array(32)(50),
      output(33) => mem_array(33)(50),
      output(34) => mem_array(34)(50),
      output(35) => mem_array(35)(50)
      );
  rom51 : entity work.rom
    generic map (
      bits  => 36,
      value => "011100000011010100000010000100010000")
    port map (
      enable_o   => mem_enable_lines(51),
      output(0)  => mem_array(0)(51),
      output(1)  => mem_array(1)(51),
      output(2)  => mem_array(2)(51),
      output(3)  => mem_array(3)(51),
      output(4)  => mem_array(4)(51),
      output(5)  => mem_array(5)(51),
      output(6)  => mem_array(6)(51),
      output(7)  => mem_array(7)(51),
      output(8)  => mem_array(8)(51),
      output(9)  => mem_array(9)(51),
      output(10) => mem_array(10)(51),
      output(11) => mem_array(11)(51),
      output(12) => mem_array(12)(51),
      output(13) => mem_array(13)(51),
      output(14) => mem_array(14)(51),
      output(15) => mem_array(15)(51),
      output(16) => mem_array(16)(51),
      output(17) => mem_array(17)(51),
      output(18) => mem_array(18)(51),
      output(19) => mem_array(19)(51),
      output(20) => mem_array(20)(51),
      output(21) => mem_array(21)(51),
      output(22) => mem_array(22)(51),
      output(23) => mem_array(23)(51),
      output(24) => mem_array(24)(51),
      output(25) => mem_array(25)(51),
      output(26) => mem_array(26)(51),
      output(27) => mem_array(27)(51),
      output(28) => mem_array(28)(51),
      output(29) => mem_array(29)(51),
      output(30) => mem_array(30)(51),
      output(31) => mem_array(31)(51),
      output(32) => mem_array(32)(51),
      output(33) => mem_array(33)(51),
      output(34) => mem_array(34)(51),
      output(35) => mem_array(35)(51)
      );
  rom52 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000010000001111000000000101000010")
    port map (
      enable_o   => mem_enable_lines(52),
      output(0)  => mem_array(0)(52),
      output(1)  => mem_array(1)(52),
      output(2)  => mem_array(2)(52),
      output(3)  => mem_array(3)(52),
      output(4)  => mem_array(4)(52),
      output(5)  => mem_array(5)(52),
      output(6)  => mem_array(6)(52),
      output(7)  => mem_array(7)(52),
      output(8)  => mem_array(8)(52),
      output(9)  => mem_array(9)(52),
      output(10) => mem_array(10)(52),
      output(11) => mem_array(11)(52),
      output(12) => mem_array(12)(52),
      output(13) => mem_array(13)(52),
      output(14) => mem_array(14)(52),
      output(15) => mem_array(15)(52),
      output(16) => mem_array(16)(52),
      output(17) => mem_array(17)(52),
      output(18) => mem_array(18)(52),
      output(19) => mem_array(19)(52),
      output(20) => mem_array(20)(52),
      output(21) => mem_array(21)(52),
      output(22) => mem_array(22)(52),
      output(23) => mem_array(23)(52),
      output(24) => mem_array(24)(52),
      output(25) => mem_array(25)(52),
      output(26) => mem_array(26)(52),
      output(27) => mem_array(27)(52),
      output(28) => mem_array(28)(52),
      output(29) => mem_array(29)(52),
      output(30) => mem_array(30)(52),
      output(31) => mem_array(31)(52),
      output(32) => mem_array(32)(52),
      output(33) => mem_array(33)(52),
      output(34) => mem_array(34)(52),
      output(35) => mem_array(35)(52)
      );
  rom53 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000011000000000110101000000100001")
    port map (
      enable_o   => mem_enable_lines(53),
      output(0)  => mem_array(0)(53),
      output(1)  => mem_array(1)(53),
      output(2)  => mem_array(2)(53),
      output(3)  => mem_array(3)(53),
      output(4)  => mem_array(4)(53),
      output(5)  => mem_array(5)(53),
      output(6)  => mem_array(6)(53),
      output(7)  => mem_array(7)(53),
      output(8)  => mem_array(8)(53),
      output(9)  => mem_array(9)(53),
      output(10) => mem_array(10)(53),
      output(11) => mem_array(11)(53),
      output(12) => mem_array(12)(53),
      output(13) => mem_array(13)(53),
      output(14) => mem_array(14)(53),
      output(15) => mem_array(15)(53),
      output(16) => mem_array(16)(53),
      output(17) => mem_array(17)(53),
      output(18) => mem_array(18)(53),
      output(19) => mem_array(19)(53),
      output(20) => mem_array(20)(53),
      output(21) => mem_array(21)(53),
      output(22) => mem_array(22)(53),
      output(23) => mem_array(23)(53),
      output(24) => mem_array(24)(53),
      output(25) => mem_array(25)(53),
      output(26) => mem_array(26)(53),
      output(27) => mem_array(27)(53),
      output(28) => mem_array(28)(53),
      output(29) => mem_array(29)(53),
      output(30) => mem_array(30)(53),
      output(31) => mem_array(31)(53),
      output(32) => mem_array(32)(53),
      output(33) => mem_array(33)(53),
      output(34) => mem_array(34)(53),
      output(35) => mem_array(35)(53)
      );
  rom54 : entity work.rom
    generic map (
      bits  => 36,
      value => "000100000001100010001001010010000000")
    port map (
      enable_o   => mem_enable_lines(54),
      output(0)  => mem_array(0)(54),
      output(1)  => mem_array(1)(54),
      output(2)  => mem_array(2)(54),
      output(3)  => mem_array(3)(54),
      output(4)  => mem_array(4)(54),
      output(5)  => mem_array(5)(54),
      output(6)  => mem_array(6)(54),
      output(7)  => mem_array(7)(54),
      output(8)  => mem_array(8)(54),
      output(9)  => mem_array(9)(54),
      output(10) => mem_array(10)(54),
      output(11) => mem_array(11)(54),
      output(12) => mem_array(12)(54),
      output(13) => mem_array(13)(54),
      output(14) => mem_array(14)(54),
      output(15) => mem_array(15)(54),
      output(16) => mem_array(16)(54),
      output(17) => mem_array(17)(54),
      output(18) => mem_array(18)(54),
      output(19) => mem_array(19)(54),
      output(20) => mem_array(20)(54),
      output(21) => mem_array(21)(54),
      output(22) => mem_array(22)(54),
      output(23) => mem_array(23)(54),
      output(24) => mem_array(24)(54),
      output(25) => mem_array(25)(54),
      output(26) => mem_array(26)(54),
      output(27) => mem_array(27)(54),
      output(28) => mem_array(28)(54),
      output(29) => mem_array(29)(54),
      output(30) => mem_array(30)(54),
      output(31) => mem_array(31)(54),
      output(32) => mem_array(32)(54),
      output(33) => mem_array(33)(54),
      output(34) => mem_array(34)(54),
      output(35) => mem_array(35)(54)
      );
  rom55 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000100000000110010000000111001000")
    port map (
      enable_o   => mem_enable_lines(55),
      output(0)  => mem_array(0)(55),
      output(1)  => mem_array(1)(55),
      output(2)  => mem_array(2)(55),
      output(3)  => mem_array(3)(55),
      output(4)  => mem_array(4)(55),
      output(5)  => mem_array(5)(55),
      output(6)  => mem_array(6)(55),
      output(7)  => mem_array(7)(55),
      output(8)  => mem_array(8)(55),
      output(9)  => mem_array(9)(55),
      output(10) => mem_array(10)(55),
      output(11) => mem_array(11)(55),
      output(12) => mem_array(12)(55),
      output(13) => mem_array(13)(55),
      output(14) => mem_array(14)(55),
      output(15) => mem_array(15)(55),
      output(16) => mem_array(16)(55),
      output(17) => mem_array(17)(55),
      output(18) => mem_array(18)(55),
      output(19) => mem_array(19)(55),
      output(20) => mem_array(20)(55),
      output(21) => mem_array(21)(55),
      output(22) => mem_array(22)(55),
      output(23) => mem_array(23)(55),
      output(24) => mem_array(24)(55),
      output(25) => mem_array(25)(55),
      output(26) => mem_array(26)(55),
      output(27) => mem_array(27)(55),
      output(28) => mem_array(28)(55),
      output(29) => mem_array(29)(55),
      output(30) => mem_array(30)(55),
      output(31) => mem_array(31)(55),
      output(32) => mem_array(32)(55),
      output(33) => mem_array(33)(55),
      output(34) => mem_array(34)(55),
      output(35) => mem_array(35)(55)
      );
  rom56 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000011000000011001100000111100")
    port map (
      enable_o   => mem_enable_lines(56),
      output(0)  => mem_array(0)(56),
      output(1)  => mem_array(1)(56),
      output(2)  => mem_array(2)(56),
      output(3)  => mem_array(3)(56),
      output(4)  => mem_array(4)(56),
      output(5)  => mem_array(5)(56),
      output(6)  => mem_array(6)(56),
      output(7)  => mem_array(7)(56),
      output(8)  => mem_array(8)(56),
      output(9)  => mem_array(9)(56),
      output(10) => mem_array(10)(56),
      output(11) => mem_array(11)(56),
      output(12) => mem_array(12)(56),
      output(13) => mem_array(13)(56),
      output(14) => mem_array(14)(56),
      output(15) => mem_array(15)(56),
      output(16) => mem_array(16)(56),
      output(17) => mem_array(17)(56),
      output(18) => mem_array(18)(56),
      output(19) => mem_array(19)(56),
      output(20) => mem_array(20)(56),
      output(21) => mem_array(21)(56),
      output(22) => mem_array(22)(56),
      output(23) => mem_array(23)(56),
      output(24) => mem_array(24)(56),
      output(25) => mem_array(25)(56),
      output(26) => mem_array(26)(56),
      output(27) => mem_array(27)(56),
      output(28) => mem_array(28)(56),
      output(29) => mem_array(29)(56),
      output(30) => mem_array(30)(56),
      output(31) => mem_array(31)(56),
      output(32) => mem_array(32)(56),
      output(33) => mem_array(33)(56),
      output(34) => mem_array(34)(56),
      output(35) => mem_array(35)(56)
      );
  rom57 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000100001100000000000000100000000")
    port map (
      enable_o   => mem_enable_lines(57),
      output(0)  => mem_array(0)(57),
      output(1)  => mem_array(1)(57),
      output(2)  => mem_array(2)(57),
      output(3)  => mem_array(3)(57),
      output(4)  => mem_array(4)(57),
      output(5)  => mem_array(5)(57),
      output(6)  => mem_array(6)(57),
      output(7)  => mem_array(7)(57),
      output(8)  => mem_array(8)(57),
      output(9)  => mem_array(9)(57),
      output(10) => mem_array(10)(57),
      output(11) => mem_array(11)(57),
      output(12) => mem_array(12)(57),
      output(13) => mem_array(13)(57),
      output(14) => mem_array(14)(57),
      output(15) => mem_array(15)(57),
      output(16) => mem_array(16)(57),
      output(17) => mem_array(17)(57),
      output(18) => mem_array(18)(57),
      output(19) => mem_array(19)(57),
      output(20) => mem_array(20)(57),
      output(21) => mem_array(21)(57),
      output(22) => mem_array(22)(57),
      output(23) => mem_array(23)(57),
      output(24) => mem_array(24)(57),
      output(25) => mem_array(25)(57),
      output(26) => mem_array(26)(57),
      output(27) => mem_array(27)(57),
      output(28) => mem_array(28)(57),
      output(29) => mem_array(29)(57),
      output(30) => mem_array(30)(57),
      output(31) => mem_array(31)(57),
      output(32) => mem_array(32)(57),
      output(33) => mem_array(33)(57),
      output(34) => mem_array(34)(57),
      output(35) => mem_array(35)(57)
      );
  rom58 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000110101000")
    port map (
      enable_o   => mem_enable_lines(58),
      output(0)  => mem_array(0)(58),
      output(1)  => mem_array(1)(58),
      output(2)  => mem_array(2)(58),
      output(3)  => mem_array(3)(58),
      output(4)  => mem_array(4)(58),
      output(5)  => mem_array(5)(58),
      output(6)  => mem_array(6)(58),
      output(7)  => mem_array(7)(58),
      output(8)  => mem_array(8)(58),
      output(9)  => mem_array(9)(58),
      output(10) => mem_array(10)(58),
      output(11) => mem_array(11)(58),
      output(12) => mem_array(12)(58),
      output(13) => mem_array(13)(58),
      output(14) => mem_array(14)(58),
      output(15) => mem_array(15)(58),
      output(16) => mem_array(16)(58),
      output(17) => mem_array(17)(58),
      output(18) => mem_array(18)(58),
      output(19) => mem_array(19)(58),
      output(20) => mem_array(20)(58),
      output(21) => mem_array(21)(58),
      output(22) => mem_array(22)(58),
      output(23) => mem_array(23)(58),
      output(24) => mem_array(24)(58),
      output(25) => mem_array(25)(58),
      output(26) => mem_array(26)(58),
      output(27) => mem_array(27)(58),
      output(28) => mem_array(28)(58),
      output(29) => mem_array(29)(58),
      output(30) => mem_array(30)(58),
      output(31) => mem_array(31)(58),
      output(32) => mem_array(32)(58),
      output(33) => mem_array(33)(58),
      output(34) => mem_array(34)(58),
      output(35) => mem_array(35)(58)
      );
  rom59 : entity work.rom
    generic map (
      bits  => 36,
      value => "000101000100000000000111000000011011")
    port map (
      enable_o   => mem_enable_lines(59),
      output(0)  => mem_array(0)(59),
      output(1)  => mem_array(1)(59),
      output(2)  => mem_array(2)(59),
      output(3)  => mem_array(3)(59),
      output(4)  => mem_array(4)(59),
      output(5)  => mem_array(5)(59),
      output(6)  => mem_array(6)(59),
      output(7)  => mem_array(7)(59),
      output(8)  => mem_array(8)(59),
      output(9)  => mem_array(9)(59),
      output(10) => mem_array(10)(59),
      output(11) => mem_array(11)(59),
      output(12) => mem_array(12)(59),
      output(13) => mem_array(13)(59),
      output(14) => mem_array(14)(59),
      output(15) => mem_array(15)(59),
      output(16) => mem_array(16)(59),
      output(17) => mem_array(17)(59),
      output(18) => mem_array(18)(59),
      output(19) => mem_array(19)(59),
      output(20) => mem_array(20)(59),
      output(21) => mem_array(21)(59),
      output(22) => mem_array(22)(59),
      output(23) => mem_array(23)(59),
      output(24) => mem_array(24)(59),
      output(25) => mem_array(25)(59),
      output(26) => mem_array(26)(59),
      output(27) => mem_array(27)(59),
      output(28) => mem_array(28)(59),
      output(29) => mem_array(29)(59),
      output(30) => mem_array(30)(59),
      output(31) => mem_array(31)(59),
      output(32) => mem_array(32)(59),
      output(33) => mem_array(33)(59),
      output(34) => mem_array(34)(59),
      output(35) => mem_array(35)(59)
      );
  rom60 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000010100001000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(60),
      output(0)  => mem_array(0)(60),
      output(1)  => mem_array(1)(60),
      output(2)  => mem_array(2)(60),
      output(3)  => mem_array(3)(60),
      output(4)  => mem_array(4)(60),
      output(5)  => mem_array(5)(60),
      output(6)  => mem_array(6)(60),
      output(7)  => mem_array(7)(60),
      output(8)  => mem_array(8)(60),
      output(9)  => mem_array(9)(60),
      output(10) => mem_array(10)(60),
      output(11) => mem_array(11)(60),
      output(12) => mem_array(12)(60),
      output(13) => mem_array(13)(60),
      output(14) => mem_array(14)(60),
      output(15) => mem_array(15)(60),
      output(16) => mem_array(16)(60),
      output(17) => mem_array(17)(60),
      output(18) => mem_array(18)(60),
      output(19) => mem_array(19)(60),
      output(20) => mem_array(20)(60),
      output(21) => mem_array(21)(60),
      output(22) => mem_array(22)(60),
      output(23) => mem_array(23)(60),
      output(24) => mem_array(24)(60),
      output(25) => mem_array(25)(60),
      output(26) => mem_array(26)(60),
      output(27) => mem_array(27)(60),
      output(28) => mem_array(28)(60),
      output(29) => mem_array(29)(60),
      output(30) => mem_array(30)(60),
      output(31) => mem_array(31)(60),
      output(32) => mem_array(32)(60),
      output(33) => mem_array(33)(60),
      output(34) => mem_array(34)(60),
      output(35) => mem_array(35)(60)
      );
  rom61 : entity work.rom
    generic map (
      bits  => 36,
      value => "111000000001010010000000000001010000")
    port map (
      enable_o   => mem_enable_lines(61),
      output(0)  => mem_array(0)(61),
      output(1)  => mem_array(1)(61),
      output(2)  => mem_array(2)(61),
      output(3)  => mem_array(3)(61),
      output(4)  => mem_array(4)(61),
      output(5)  => mem_array(5)(61),
      output(6)  => mem_array(6)(61),
      output(7)  => mem_array(7)(61),
      output(8)  => mem_array(8)(61),
      output(9)  => mem_array(9)(61),
      output(10) => mem_array(10)(61),
      output(11) => mem_array(11)(61),
      output(12) => mem_array(12)(61),
      output(13) => mem_array(13)(61),
      output(14) => mem_array(14)(61),
      output(15) => mem_array(15)(61),
      output(16) => mem_array(16)(61),
      output(17) => mem_array(17)(61),
      output(18) => mem_array(18)(61),
      output(19) => mem_array(19)(61),
      output(20) => mem_array(20)(61),
      output(21) => mem_array(21)(61),
      output(22) => mem_array(22)(61),
      output(23) => mem_array(23)(61),
      output(24) => mem_array(24)(61),
      output(25) => mem_array(25)(61),
      output(26) => mem_array(26)(61),
      output(27) => mem_array(27)(61),
      output(28) => mem_array(28)(61),
      output(29) => mem_array(29)(61),
      output(30) => mem_array(30)(61),
      output(31) => mem_array(31)(61),
      output(32) => mem_array(32)(61),
      output(33) => mem_array(33)(61),
      output(34) => mem_array(34)(61),
      output(35) => mem_array(35)(61)
      );
  rom62 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001010000101000000000000001000")
    port map (
      enable_o   => mem_enable_lines(62),
      output(0)  => mem_array(0)(62),
      output(1)  => mem_array(1)(62),
      output(2)  => mem_array(2)(62),
      output(3)  => mem_array(3)(62),
      output(4)  => mem_array(4)(62),
      output(5)  => mem_array(5)(62),
      output(6)  => mem_array(6)(62),
      output(7)  => mem_array(7)(62),
      output(8)  => mem_array(8)(62),
      output(9)  => mem_array(9)(62),
      output(10) => mem_array(10)(62),
      output(11) => mem_array(11)(62),
      output(12) => mem_array(12)(62),
      output(13) => mem_array(13)(62),
      output(14) => mem_array(14)(62),
      output(15) => mem_array(15)(62),
      output(16) => mem_array(16)(62),
      output(17) => mem_array(17)(62),
      output(18) => mem_array(18)(62),
      output(19) => mem_array(19)(62),
      output(20) => mem_array(20)(62),
      output(21) => mem_array(21)(62),
      output(22) => mem_array(22)(62),
      output(23) => mem_array(23)(62),
      output(24) => mem_array(24)(62),
      output(25) => mem_array(25)(62),
      output(26) => mem_array(26)(62),
      output(27) => mem_array(27)(62),
      output(28) => mem_array(28)(62),
      output(29) => mem_array(29)(62),
      output(30) => mem_array(30)(62),
      output(31) => mem_array(31)(62),
      output(32) => mem_array(32)(62),
      output(33) => mem_array(33)(62),
      output(34) => mem_array(34)(62),
      output(35) => mem_array(35)(62)
      );
  rom63 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000011100100000010100010000000000")
    port map (
      enable_o   => mem_enable_lines(63),
      output(0)  => mem_array(0)(63),
      output(1)  => mem_array(1)(63),
      output(2)  => mem_array(2)(63),
      output(3)  => mem_array(3)(63),
      output(4)  => mem_array(4)(63),
      output(5)  => mem_array(5)(63),
      output(6)  => mem_array(6)(63),
      output(7)  => mem_array(7)(63),
      output(8)  => mem_array(8)(63),
      output(9)  => mem_array(9)(63),
      output(10) => mem_array(10)(63),
      output(11) => mem_array(11)(63),
      output(12) => mem_array(12)(63),
      output(13) => mem_array(13)(63),
      output(14) => mem_array(14)(63),
      output(15) => mem_array(15)(63),
      output(16) => mem_array(16)(63),
      output(17) => mem_array(17)(63),
      output(18) => mem_array(18)(63),
      output(19) => mem_array(19)(63),
      output(20) => mem_array(20)(63),
      output(21) => mem_array(21)(63),
      output(22) => mem_array(22)(63),
      output(23) => mem_array(23)(63),
      output(24) => mem_array(24)(63),
      output(25) => mem_array(25)(63),
      output(26) => mem_array(26)(63),
      output(27) => mem_array(27)(63),
      output(28) => mem_array(28)(63),
      output(29) => mem_array(29)(63),
      output(30) => mem_array(30)(63),
      output(31) => mem_array(31)(63),
      output(32) => mem_array(32)(63),
      output(33) => mem_array(33)(63),
      output(34) => mem_array(34)(63),
      output(35) => mem_array(35)(63)
      );
  rom64 : entity work.rom
    generic map (
      bits  => 36,
      value => "011100000001110100000001010000100000")
    port map (
      enable_o   => mem_enable_lines(64),
      output(0)  => mem_array(0)(64),
      output(1)  => mem_array(1)(64),
      output(2)  => mem_array(2)(64),
      output(3)  => mem_array(3)(64),
      output(4)  => mem_array(4)(64),
      output(5)  => mem_array(5)(64),
      output(6)  => mem_array(6)(64),
      output(7)  => mem_array(7)(64),
      output(8)  => mem_array(8)(64),
      output(9)  => mem_array(9)(64),
      output(10) => mem_array(10)(64),
      output(11) => mem_array(11)(64),
      output(12) => mem_array(12)(64),
      output(13) => mem_array(13)(64),
      output(14) => mem_array(14)(64),
      output(15) => mem_array(15)(64),
      output(16) => mem_array(16)(64),
      output(17) => mem_array(17)(64),
      output(18) => mem_array(18)(64),
      output(19) => mem_array(19)(64),
      output(20) => mem_array(20)(64),
      output(21) => mem_array(21)(64),
      output(22) => mem_array(22)(64),
      output(23) => mem_array(23)(64),
      output(24) => mem_array(24)(64),
      output(25) => mem_array(25)(64),
      output(26) => mem_array(26)(64),
      output(27) => mem_array(27)(64),
      output(28) => mem_array(28)(64),
      output(29) => mem_array(29)(64),
      output(30) => mem_array(30)(64),
      output(31) => mem_array(31)(64),
      output(32) => mem_array(32)(64),
      output(33) => mem_array(33)(64),
      output(34) => mem_array(34)(64),
      output(35) => mem_array(35)(64)
      );
  rom65 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000001001000101000000")
    port map (
      enable_o   => mem_enable_lines(65),
      output(0)  => mem_array(0)(65),
      output(1)  => mem_array(1)(65),
      output(2)  => mem_array(2)(65),
      output(3)  => mem_array(3)(65),
      output(4)  => mem_array(4)(65),
      output(5)  => mem_array(5)(65),
      output(6)  => mem_array(6)(65),
      output(7)  => mem_array(7)(65),
      output(8)  => mem_array(8)(65),
      output(9)  => mem_array(9)(65),
      output(10) => mem_array(10)(65),
      output(11) => mem_array(11)(65),
      output(12) => mem_array(12)(65),
      output(13) => mem_array(13)(65),
      output(14) => mem_array(14)(65),
      output(15) => mem_array(15)(65),
      output(16) => mem_array(16)(65),
      output(17) => mem_array(17)(65),
      output(18) => mem_array(18)(65),
      output(19) => mem_array(19)(65),
      output(20) => mem_array(20)(65),
      output(21) => mem_array(21)(65),
      output(22) => mem_array(22)(65),
      output(23) => mem_array(23)(65),
      output(24) => mem_array(24)(65),
      output(25) => mem_array(25)(65),
      output(26) => mem_array(26)(65),
      output(27) => mem_array(27)(65),
      output(28) => mem_array(28)(65),
      output(29) => mem_array(29)(65),
      output(30) => mem_array(30)(65),
      output(31) => mem_array(31)(65),
      output(32) => mem_array(32)(65),
      output(33) => mem_array(33)(65),
      output(34) => mem_array(34)(65),
      output(35) => mem_array(35)(65)
      );
  rom66 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001000000000011110000000110110")
    port map (
      enable_o   => mem_enable_lines(66),
      output(0)  => mem_array(0)(66),
      output(1)  => mem_array(1)(66),
      output(2)  => mem_array(2)(66),
      output(3)  => mem_array(3)(66),
      output(4)  => mem_array(4)(66),
      output(5)  => mem_array(5)(66),
      output(6)  => mem_array(6)(66),
      output(7)  => mem_array(7)(66),
      output(8)  => mem_array(8)(66),
      output(9)  => mem_array(9)(66),
      output(10) => mem_array(10)(66),
      output(11) => mem_array(11)(66),
      output(12) => mem_array(12)(66),
      output(13) => mem_array(13)(66),
      output(14) => mem_array(14)(66),
      output(15) => mem_array(15)(66),
      output(16) => mem_array(16)(66),
      output(17) => mem_array(17)(66),
      output(18) => mem_array(18)(66),
      output(19) => mem_array(19)(66),
      output(20) => mem_array(20)(66),
      output(21) => mem_array(21)(66),
      output(22) => mem_array(22)(66),
      output(23) => mem_array(23)(66),
      output(24) => mem_array(24)(66),
      output(25) => mem_array(25)(66),
      output(26) => mem_array(26)(66),
      output(27) => mem_array(27)(66),
      output(28) => mem_array(28)(66),
      output(29) => mem_array(29)(66),
      output(30) => mem_array(30)(66),
      output(31) => mem_array(31)(66),
      output(32) => mem_array(32)(66),
      output(33) => mem_array(33)(66),
      output(34) => mem_array(34)(66),
      output(35) => mem_array(35)(66)
      );
  rom67 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001001000010000000001111010000001")
    port map (
      enable_o   => mem_enable_lines(67),
      output(0)  => mem_array(0)(67),
      output(1)  => mem_array(1)(67),
      output(2)  => mem_array(2)(67),
      output(3)  => mem_array(3)(67),
      output(4)  => mem_array(4)(67),
      output(5)  => mem_array(5)(67),
      output(6)  => mem_array(6)(67),
      output(7)  => mem_array(7)(67),
      output(8)  => mem_array(8)(67),
      output(9)  => mem_array(9)(67),
      output(10) => mem_array(10)(67),
      output(11) => mem_array(11)(67),
      output(12) => mem_array(12)(67),
      output(13) => mem_array(13)(67),
      output(14) => mem_array(14)(67),
      output(15) => mem_array(15)(67),
      output(16) => mem_array(16)(67),
      output(17) => mem_array(17)(67),
      output(18) => mem_array(18)(67),
      output(19) => mem_array(19)(67),
      output(20) => mem_array(20)(67),
      output(21) => mem_array(21)(67),
      output(22) => mem_array(22)(67),
      output(23) => mem_array(23)(67),
      output(24) => mem_array(24)(67),
      output(25) => mem_array(25)(67),
      output(26) => mem_array(26)(67),
      output(27) => mem_array(27)(67),
      output(28) => mem_array(28)(67),
      output(29) => mem_array(29)(67),
      output(30) => mem_array(30)(67),
      output(31) => mem_array(31)(67),
      output(32) => mem_array(32)(67),
      output(33) => mem_array(33)(67),
      output(34) => mem_array(34)(67),
      output(35) => mem_array(35)(67)
      );
  rom68 : entity work.rom
    generic map (
      bits  => 36,
      value => "010010000000001000000000000111110000")
    port map (
      enable_o   => mem_enable_lines(68),
      output(0)  => mem_array(0)(68),
      output(1)  => mem_array(1)(68),
      output(2)  => mem_array(2)(68),
      output(3)  => mem_array(3)(68),
      output(4)  => mem_array(4)(68),
      output(5)  => mem_array(5)(68),
      output(6)  => mem_array(6)(68),
      output(7)  => mem_array(7)(68),
      output(8)  => mem_array(8)(68),
      output(9)  => mem_array(9)(68),
      output(10) => mem_array(10)(68),
      output(11) => mem_array(11)(68),
      output(12) => mem_array(12)(68),
      output(13) => mem_array(13)(68),
      output(14) => mem_array(14)(68),
      output(15) => mem_array(15)(68),
      output(16) => mem_array(16)(68),
      output(17) => mem_array(17)(68),
      output(18) => mem_array(18)(68),
      output(19) => mem_array(19)(68),
      output(20) => mem_array(20)(68),
      output(21) => mem_array(21)(68),
      output(22) => mem_array(22)(68),
      output(23) => mem_array(23)(68),
      output(24) => mem_array(24)(68),
      output(25) => mem_array(25)(68),
      output(26) => mem_array(26)(68),
      output(27) => mem_array(27)(68),
      output(28) => mem_array(28)(68),
      output(29) => mem_array(29)(68),
      output(30) => mem_array(30)(68),
      output(31) => mem_array(31)(68),
      output(32) => mem_array(32)(68),
      output(33) => mem_array(33)(68),
      output(34) => mem_array(34)(68),
      output(35) => mem_array(35)(68)
      );
  rom69 : entity work.rom
    generic map (
      bits  => 36,
      value => "000101000100000000000111000000011111")
    port map (
      enable_o   => mem_enable_lines(69),
      output(0)  => mem_array(0)(69),
      output(1)  => mem_array(1)(69),
      output(2)  => mem_array(2)(69),
      output(3)  => mem_array(3)(69),
      output(4)  => mem_array(4)(69),
      output(5)  => mem_array(5)(69),
      output(6)  => mem_array(6)(69),
      output(7)  => mem_array(7)(69),
      output(8)  => mem_array(8)(69),
      output(9)  => mem_array(9)(69),
      output(10) => mem_array(10)(69),
      output(11) => mem_array(11)(69),
      output(12) => mem_array(12)(69),
      output(13) => mem_array(13)(69),
      output(14) => mem_array(14)(69),
      output(15) => mem_array(15)(69),
      output(16) => mem_array(16)(69),
      output(17) => mem_array(17)(69),
      output(18) => mem_array(18)(69),
      output(19) => mem_array(19)(69),
      output(20) => mem_array(20)(69),
      output(21) => mem_array(21)(69),
      output(22) => mem_array(22)(69),
      output(23) => mem_array(23)(69),
      output(24) => mem_array(24)(69),
      output(25) => mem_array(25)(69),
      output(26) => mem_array(26)(69),
      output(27) => mem_array(27)(69),
      output(28) => mem_array(28)(69),
      output(29) => mem_array(29)(69),
      output(30) => mem_array(30)(69),
      output(31) => mem_array(31)(69),
      output(32) => mem_array(32)(69),
      output(33) => mem_array(33)(69),
      output(34) => mem_array(34)(69),
      output(35) => mem_array(35)(69)
      );
  rom70 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000010100001000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(70),
      output(0)  => mem_array(0)(70),
      output(1)  => mem_array(1)(70),
      output(2)  => mem_array(2)(70),
      output(3)  => mem_array(3)(70),
      output(4)  => mem_array(4)(70),
      output(5)  => mem_array(5)(70),
      output(6)  => mem_array(6)(70),
      output(7)  => mem_array(7)(70),
      output(8)  => mem_array(8)(70),
      output(9)  => mem_array(9)(70),
      output(10) => mem_array(10)(70),
      output(11) => mem_array(11)(70),
      output(12) => mem_array(12)(70),
      output(13) => mem_array(13)(70),
      output(14) => mem_array(14)(70),
      output(15) => mem_array(15)(70),
      output(16) => mem_array(16)(70),
      output(17) => mem_array(17)(70),
      output(18) => mem_array(18)(70),
      output(19) => mem_array(19)(70),
      output(20) => mem_array(20)(70),
      output(21) => mem_array(21)(70),
      output(22) => mem_array(22)(70),
      output(23) => mem_array(23)(70),
      output(24) => mem_array(24)(70),
      output(25) => mem_array(25)(70),
      output(26) => mem_array(26)(70),
      output(27) => mem_array(27)(70),
      output(28) => mem_array(28)(70),
      output(29) => mem_array(29)(70),
      output(30) => mem_array(30)(70),
      output(31) => mem_array(31)(70),
      output(32) => mem_array(32)(70),
      output(33) => mem_array(33)(70),
      output(34) => mem_array(34)(70),
      output(35) => mem_array(35)(70)
      );
  rom71 : entity work.rom
    generic map (
      bits  => 36,
      value => "000010010011111100000000000010000000")
    port map (
      enable_o   => mem_enable_lines(71),
      output(0)  => mem_array(0)(71),
      output(1)  => mem_array(1)(71),
      output(2)  => mem_array(2)(71),
      output(3)  => mem_array(3)(71),
      output(4)  => mem_array(4)(71),
      output(5)  => mem_array(5)(71),
      output(6)  => mem_array(6)(71),
      output(7)  => mem_array(7)(71),
      output(8)  => mem_array(8)(71),
      output(9)  => mem_array(9)(71),
      output(10) => mem_array(10)(71),
      output(11) => mem_array(11)(71),
      output(12) => mem_array(12)(71),
      output(13) => mem_array(13)(71),
      output(14) => mem_array(14)(71),
      output(15) => mem_array(15)(71),
      output(16) => mem_array(16)(71),
      output(17) => mem_array(17)(71),
      output(18) => mem_array(18)(71),
      output(19) => mem_array(19)(71),
      output(20) => mem_array(20)(71),
      output(21) => mem_array(21)(71),
      output(22) => mem_array(22)(71),
      output(23) => mem_array(23)(71),
      output(24) => mem_array(24)(71),
      output(25) => mem_array(25)(71),
      output(26) => mem_array(26)(71),
      output(27) => mem_array(27)(71),
      output(28) => mem_array(28)(71),
      output(29) => mem_array(29)(71),
      output(30) => mem_array(30)(71),
      output(31) => mem_array(31)(71),
      output(32) => mem_array(32)(71),
      output(33) => mem_array(33)(71),
      output(34) => mem_array(34)(71),
      output(35) => mem_array(35)(71)
      );
  rom72 : entity work.rom
    generic map (
      bits  => 36,
      value => "001000001000001101010000001000010001")
    port map (
      enable_o   => mem_enable_lines(72),
      output(0)  => mem_array(0)(72),
      output(1)  => mem_array(1)(72),
      output(2)  => mem_array(2)(72),
      output(3)  => mem_array(3)(72),
      output(4)  => mem_array(4)(72),
      output(5)  => mem_array(5)(72),
      output(6)  => mem_array(6)(72),
      output(7)  => mem_array(7)(72),
      output(8)  => mem_array(8)(72),
      output(9)  => mem_array(9)(72),
      output(10) => mem_array(10)(72),
      output(11) => mem_array(11)(72),
      output(12) => mem_array(12)(72),
      output(13) => mem_array(13)(72),
      output(14) => mem_array(14)(72),
      output(15) => mem_array(15)(72),
      output(16) => mem_array(16)(72),
      output(17) => mem_array(17)(72),
      output(18) => mem_array(18)(72),
      output(19) => mem_array(19)(72),
      output(20) => mem_array(20)(72),
      output(21) => mem_array(21)(72),
      output(22) => mem_array(22)(72),
      output(23) => mem_array(23)(72),
      output(24) => mem_array(24)(72),
      output(25) => mem_array(25)(72),
      output(26) => mem_array(26)(72),
      output(27) => mem_array(27)(72),
      output(28) => mem_array(28)(72),
      output(29) => mem_array(29)(72),
      output(30) => mem_array(30)(72),
      output(31) => mem_array(31)(72),
      output(32) => mem_array(32)(72),
      output(33) => mem_array(33)(72),
      output(34) => mem_array(34)(72),
      output(35) => mem_array(35)(72)
      );
  rom73 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000001000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(73),
      output(0)  => mem_array(0)(73),
      output(1)  => mem_array(1)(73),
      output(2)  => mem_array(2)(73),
      output(3)  => mem_array(3)(73),
      output(4)  => mem_array(4)(73),
      output(5)  => mem_array(5)(73),
      output(6)  => mem_array(6)(73),
      output(7)  => mem_array(7)(73),
      output(8)  => mem_array(8)(73),
      output(9)  => mem_array(9)(73),
      output(10) => mem_array(10)(73),
      output(11) => mem_array(11)(73),
      output(12) => mem_array(12)(73),
      output(13) => mem_array(13)(73),
      output(14) => mem_array(14)(73),
      output(15) => mem_array(15)(73),
      output(16) => mem_array(16)(73),
      output(17) => mem_array(17)(73),
      output(18) => mem_array(18)(73),
      output(19) => mem_array(19)(73),
      output(20) => mem_array(20)(73),
      output(21) => mem_array(21)(73),
      output(22) => mem_array(22)(73),
      output(23) => mem_array(23)(73),
      output(24) => mem_array(24)(73),
      output(25) => mem_array(25)(73),
      output(26) => mem_array(26)(73),
      output(27) => mem_array(27)(73),
      output(28) => mem_array(28)(73),
      output(29) => mem_array(29)(73),
      output(30) => mem_array(30)(73),
      output(31) => mem_array(31)(73),
      output(32) => mem_array(32)(73),
      output(33) => mem_array(33)(73),
      output(34) => mem_array(34)(73),
      output(35) => mem_array(35)(73)
      );
  rom74 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000010000110001001010010000000")
    port map (
      enable_o   => mem_enable_lines(74),
      output(0)  => mem_array(0)(74),
      output(1)  => mem_array(1)(74),
      output(2)  => mem_array(2)(74),
      output(3)  => mem_array(3)(74),
      output(4)  => mem_array(4)(74),
      output(5)  => mem_array(5)(74),
      output(6)  => mem_array(6)(74),
      output(7)  => mem_array(7)(74),
      output(8)  => mem_array(8)(74),
      output(9)  => mem_array(9)(74),
      output(10) => mem_array(10)(74),
      output(11) => mem_array(11)(74),
      output(12) => mem_array(12)(74),
      output(13) => mem_array(13)(74),
      output(14) => mem_array(14)(74),
      output(15) => mem_array(15)(74),
      output(16) => mem_array(16)(74),
      output(17) => mem_array(17)(74),
      output(18) => mem_array(18)(74),
      output(19) => mem_array(19)(74),
      output(20) => mem_array(20)(74),
      output(21) => mem_array(21)(74),
      output(22) => mem_array(22)(74),
      output(23) => mem_array(23)(74),
      output(24) => mem_array(24)(74),
      output(25) => mem_array(25)(74),
      output(26) => mem_array(26)(74),
      output(27) => mem_array(27)(74),
      output(28) => mem_array(28)(74),
      output(29) => mem_array(29)(74),
      output(30) => mem_array(30)(74),
      output(31) => mem_array(31)(74),
      output(32) => mem_array(32)(74),
      output(33) => mem_array(33)(74),
      output(34) => mem_array(34)(74),
      output(35) => mem_array(35)(74)
      );
  rom75 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000110000001000100000000111001000")
    port map (
      enable_o   => mem_enable_lines(75),
      output(0)  => mem_array(0)(75),
      output(1)  => mem_array(1)(75),
      output(2)  => mem_array(2)(75),
      output(3)  => mem_array(3)(75),
      output(4)  => mem_array(4)(75),
      output(5)  => mem_array(5)(75),
      output(6)  => mem_array(6)(75),
      output(7)  => mem_array(7)(75),
      output(8)  => mem_array(8)(75),
      output(9)  => mem_array(9)(75),
      output(10) => mem_array(10)(75),
      output(11) => mem_array(11)(75),
      output(12) => mem_array(12)(75),
      output(13) => mem_array(13)(75),
      output(14) => mem_array(14)(75),
      output(15) => mem_array(15)(75),
      output(16) => mem_array(16)(75),
      output(17) => mem_array(17)(75),
      output(18) => mem_array(18)(75),
      output(19) => mem_array(19)(75),
      output(20) => mem_array(20)(75),
      output(21) => mem_array(21)(75),
      output(22) => mem_array(22)(75),
      output(23) => mem_array(23)(75),
      output(24) => mem_array(24)(75),
      output(25) => mem_array(25)(75),
      output(26) => mem_array(26)(75),
      output(27) => mem_array(27)(75),
      output(28) => mem_array(28)(75),
      output(29) => mem_array(29)(75),
      output(30) => mem_array(30)(75),
      output(31) => mem_array(31)(75),
      output(32) => mem_array(32)(75),
      output(33) => mem_array(33)(75),
      output(34) => mem_array(34)(75),
      output(35) => mem_array(35)(75)
      );
  rom76 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000011000000100010100000111100")
    port map (
      enable_o   => mem_enable_lines(76),
      output(0)  => mem_array(0)(76),
      output(1)  => mem_array(1)(76),
      output(2)  => mem_array(2)(76),
      output(3)  => mem_array(3)(76),
      output(4)  => mem_array(4)(76),
      output(5)  => mem_array(5)(76),
      output(6)  => mem_array(6)(76),
      output(7)  => mem_array(7)(76),
      output(8)  => mem_array(8)(76),
      output(9)  => mem_array(9)(76),
      output(10) => mem_array(10)(76),
      output(11) => mem_array(11)(76),
      output(12) => mem_array(12)(76),
      output(13) => mem_array(13)(76),
      output(14) => mem_array(14)(76),
      output(15) => mem_array(15)(76),
      output(16) => mem_array(16)(76),
      output(17) => mem_array(17)(76),
      output(18) => mem_array(18)(76),
      output(19) => mem_array(19)(76),
      output(20) => mem_array(20)(76),
      output(21) => mem_array(21)(76),
      output(22) => mem_array(22)(76),
      output(23) => mem_array(23)(76),
      output(24) => mem_array(24)(76),
      output(25) => mem_array(25)(76),
      output(26) => mem_array(26)(76),
      output(27) => mem_array(27)(76),
      output(28) => mem_array(28)(76),
      output(29) => mem_array(29)(76),
      output(30) => mem_array(30)(76),
      output(31) => mem_array(31)(76),
      output(32) => mem_array(32)(76),
      output(33) => mem_array(33)(76),
      output(34) => mem_array(34)(76),
      output(35) => mem_array(35)(76)
      );
  rom77 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001010011000000010001100000011")
    port map (
      enable_o   => mem_enable_lines(77),
      output(0)  => mem_array(0)(77),
      output(1)  => mem_array(1)(77),
      output(2)  => mem_array(2)(77),
      output(3)  => mem_array(3)(77),
      output(4)  => mem_array(4)(77),
      output(5)  => mem_array(5)(77),
      output(6)  => mem_array(6)(77),
      output(7)  => mem_array(7)(77),
      output(8)  => mem_array(8)(77),
      output(9)  => mem_array(9)(77),
      output(10) => mem_array(10)(77),
      output(11) => mem_array(11)(77),
      output(12) => mem_array(12)(77),
      output(13) => mem_array(13)(77),
      output(14) => mem_array(14)(77),
      output(15) => mem_array(15)(77),
      output(16) => mem_array(16)(77),
      output(17) => mem_array(17)(77),
      output(18) => mem_array(18)(77),
      output(19) => mem_array(19)(77),
      output(20) => mem_array(20)(77),
      output(21) => mem_array(21)(77),
      output(22) => mem_array(22)(77),
      output(23) => mem_array(23)(77),
      output(24) => mem_array(24)(77),
      output(25) => mem_array(25)(77),
      output(26) => mem_array(26)(77),
      output(27) => mem_array(27)(77),
      output(28) => mem_array(28)(77),
      output(29) => mem_array(29)(77),
      output(30) => mem_array(30)(77),
      output(31) => mem_array(31)(77),
      output(32) => mem_array(32)(77),
      output(33) => mem_array(33)(77),
      output(34) => mem_array(34)(77),
      output(35) => mem_array(35)(77)
      );
  rom78 : entity work.rom
    generic map (
      bits  => 36,
      value => "010101000000000000010000001000111000")
    port map (
      enable_o   => mem_enable_lines(78),
      output(0)  => mem_array(0)(78),
      output(1)  => mem_array(1)(78),
      output(2)  => mem_array(2)(78),
      output(3)  => mem_array(3)(78),
      output(4)  => mem_array(4)(78),
      output(5)  => mem_array(5)(78),
      output(6)  => mem_array(6)(78),
      output(7)  => mem_array(7)(78),
      output(8)  => mem_array(8)(78),
      output(9)  => mem_array(9)(78),
      output(10) => mem_array(10)(78),
      output(11) => mem_array(11)(78),
      output(12) => mem_array(12)(78),
      output(13) => mem_array(13)(78),
      output(14) => mem_array(14)(78),
      output(15) => mem_array(15)(78),
      output(16) => mem_array(16)(78),
      output(17) => mem_array(17)(78),
      output(18) => mem_array(18)(78),
      output(19) => mem_array(19)(78),
      output(20) => mem_array(20)(78),
      output(21) => mem_array(21)(78),
      output(22) => mem_array(22)(78),
      output(23) => mem_array(23)(78),
      output(24) => mem_array(24)(78),
      output(25) => mem_array(25)(78),
      output(26) => mem_array(26)(78),
      output(27) => mem_array(27)(78),
      output(28) => mem_array(28)(78),
      output(29) => mem_array(29)(78),
      output(30) => mem_array(30)(78),
      output(31) => mem_array(31)(78),
      output(32) => mem_array(32)(78),
      output(33) => mem_array(33)(78),
      output(34) => mem_array(34)(78),
      output(35) => mem_array(35)(78)
      );
  rom79 : entity work.rom
    generic map (
      bits  => 36,
      value => "000101000000001000010000000000100100")
    port map (
      enable_o   => mem_enable_lines(79),
      output(0)  => mem_array(0)(79),
      output(1)  => mem_array(1)(79),
      output(2)  => mem_array(2)(79),
      output(3)  => mem_array(3)(79),
      output(4)  => mem_array(4)(79),
      output(5)  => mem_array(5)(79),
      output(6)  => mem_array(6)(79),
      output(7)  => mem_array(7)(79),
      output(8)  => mem_array(8)(79),
      output(9)  => mem_array(9)(79),
      output(10) => mem_array(10)(79),
      output(11) => mem_array(11)(79),
      output(12) => mem_array(12)(79),
      output(13) => mem_array(13)(79),
      output(14) => mem_array(14)(79),
      output(15) => mem_array(15)(79),
      output(16) => mem_array(16)(79),
      output(17) => mem_array(17)(79),
      output(18) => mem_array(18)(79),
      output(19) => mem_array(19)(79),
      output(20) => mem_array(20)(79),
      output(21) => mem_array(21)(79),
      output(22) => mem_array(22)(79),
      output(23) => mem_array(23)(79),
      output(24) => mem_array(24)(79),
      output(25) => mem_array(25)(79),
      output(26) => mem_array(26)(79),
      output(27) => mem_array(27)(79),
      output(28) => mem_array(28)(79),
      output(29) => mem_array(29)(79),
      output(30) => mem_array(30)(79),
      output(31) => mem_array(31)(79),
      output(32) => mem_array(32)(79),
      output(33) => mem_array(33)(79),
      output(34) => mem_array(34)(79),
      output(35) => mem_array(35)(79)
      );
  rom80 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000110101000000100001000100000010")
    port map (
      enable_o   => mem_enable_lines(80),
      output(0)  => mem_array(0)(80),
      output(1)  => mem_array(1)(80),
      output(2)  => mem_array(2)(80),
      output(3)  => mem_array(3)(80),
      output(4)  => mem_array(4)(80),
      output(5)  => mem_array(5)(80),
      output(6)  => mem_array(6)(80),
      output(7)  => mem_array(7)(80),
      output(8)  => mem_array(8)(80),
      output(9)  => mem_array(9)(80),
      output(10) => mem_array(10)(80),
      output(11) => mem_array(11)(80),
      output(12) => mem_array(12)(80),
      output(13) => mem_array(13)(80),
      output(14) => mem_array(14)(80),
      output(15) => mem_array(15)(80),
      output(16) => mem_array(16)(80),
      output(17) => mem_array(17)(80),
      output(18) => mem_array(18)(80),
      output(19) => mem_array(19)(80),
      output(20) => mem_array(20)(80),
      output(21) => mem_array(21)(80),
      output(22) => mem_array(22)(80),
      output(23) => mem_array(23)(80),
      output(24) => mem_array(24)(80),
      output(25) => mem_array(25)(80),
      output(26) => mem_array(26)(80),
      output(27) => mem_array(27)(80),
      output(28) => mem_array(28)(80),
      output(29) => mem_array(29)(80),
      output(30) => mem_array(30)(80),
      output(31) => mem_array(31)(80),
      output(32) => mem_array(32)(80),
      output(33) => mem_array(33)(80),
      output(34) => mem_array(34)(80),
      output(35) => mem_array(35)(80)
      );
  rom81 : entity work.rom
    generic map (
      bits  => 36,
      value => "010010001001010010000000000000110000")
    port map (
      enable_o   => mem_enable_lines(81),
      output(0)  => mem_array(0)(81),
      output(1)  => mem_array(1)(81),
      output(2)  => mem_array(2)(81),
      output(3)  => mem_array(3)(81),
      output(4)  => mem_array(4)(81),
      output(5)  => mem_array(5)(81),
      output(6)  => mem_array(6)(81),
      output(7)  => mem_array(7)(81),
      output(8)  => mem_array(8)(81),
      output(9)  => mem_array(9)(81),
      output(10) => mem_array(10)(81),
      output(11) => mem_array(11)(81),
      output(12) => mem_array(12)(81),
      output(13) => mem_array(13)(81),
      output(14) => mem_array(14)(81),
      output(15) => mem_array(15)(81),
      output(16) => mem_array(16)(81),
      output(17) => mem_array(17)(81),
      output(18) => mem_array(18)(81),
      output(19) => mem_array(19)(81),
      output(20) => mem_array(20)(81),
      output(21) => mem_array(21)(81),
      output(22) => mem_array(22)(81),
      output(23) => mem_array(23)(81),
      output(24) => mem_array(24)(81),
      output(25) => mem_array(25)(81),
      output(26) => mem_array(26)(81),
      output(27) => mem_array(27)(81),
      output(28) => mem_array(28)(81),
      output(29) => mem_array(29)(81),
      output(30) => mem_array(30)(81),
      output(31) => mem_array(31)(81),
      output(32) => mem_array(32)(81),
      output(33) => mem_array(33)(81),
      output(34) => mem_array(34)(81),
      output(35) => mem_array(35)(81)
      );
  rom82 : entity work.rom
    generic map (
      bits  => 36,
      value => "001001010000000111001000000000000011")
    port map (
      enable_o   => mem_enable_lines(82),
      output(0)  => mem_array(0)(82),
      output(1)  => mem_array(1)(82),
      output(2)  => mem_array(2)(82),
      output(3)  => mem_array(3)(82),
      output(4)  => mem_array(4)(82),
      output(5)  => mem_array(5)(82),
      output(6)  => mem_array(6)(82),
      output(7)  => mem_array(7)(82),
      output(8)  => mem_array(8)(82),
      output(9)  => mem_array(9)(82),
      output(10) => mem_array(10)(82),
      output(11) => mem_array(11)(82),
      output(12) => mem_array(12)(82),
      output(13) => mem_array(13)(82),
      output(14) => mem_array(14)(82),
      output(15) => mem_array(15)(82),
      output(16) => mem_array(16)(82),
      output(17) => mem_array(17)(82),
      output(18) => mem_array(18)(82),
      output(19) => mem_array(19)(82),
      output(20) => mem_array(20)(82),
      output(21) => mem_array(21)(82),
      output(22) => mem_array(22)(82),
      output(23) => mem_array(23)(82),
      output(24) => mem_array(24)(82),
      output(25) => mem_array(25)(82),
      output(26) => mem_array(26)(82),
      output(27) => mem_array(27)(82),
      output(28) => mem_array(28)(82),
      output(29) => mem_array(29)(82),
      output(30) => mem_array(30)(82),
      output(31) => mem_array(31)(82),
      output(32) => mem_array(32)(82),
      output(33) => mem_array(33)(82),
      output(34) => mem_array(34)(82),
      output(35) => mem_array(35)(82)
      );
  rom83 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000100101100000110101000000100001")
    port map (
      enable_o   => mem_enable_lines(83),
      output(0)  => mem_array(0)(83),
      output(1)  => mem_array(1)(83),
      output(2)  => mem_array(2)(83),
      output(3)  => mem_array(3)(83),
      output(4)  => mem_array(4)(83),
      output(5)  => mem_array(5)(83),
      output(6)  => mem_array(6)(83),
      output(7)  => mem_array(7)(83),
      output(8)  => mem_array(8)(83),
      output(9)  => mem_array(9)(83),
      output(10) => mem_array(10)(83),
      output(11) => mem_array(11)(83),
      output(12) => mem_array(12)(83),
      output(13) => mem_array(13)(83),
      output(14) => mem_array(14)(83),
      output(15) => mem_array(15)(83),
      output(16) => mem_array(16)(83),
      output(17) => mem_array(17)(83),
      output(18) => mem_array(18)(83),
      output(19) => mem_array(19)(83),
      output(20) => mem_array(20)(83),
      output(21) => mem_array(21)(83),
      output(22) => mem_array(22)(83),
      output(23) => mem_array(23)(83),
      output(24) => mem_array(24)(83),
      output(25) => mem_array(25)(83),
      output(26) => mem_array(26)(83),
      output(27) => mem_array(27)(83),
      output(28) => mem_array(28)(83),
      output(29) => mem_array(29)(83),
      output(30) => mem_array(30)(83),
      output(31) => mem_array(31)(83),
      output(32) => mem_array(32)(83),
      output(33) => mem_array(33)(83),
      output(34) => mem_array(34)(83),
      output(35) => mem_array(35)(83)
      );
  rom84 : entity work.rom
    generic map (
      bits  => 36,
      value => "000100000010011000000011111100100000")
    port map (
      enable_o   => mem_enable_lines(84),
      output(0)  => mem_array(0)(84),
      output(1)  => mem_array(1)(84),
      output(2)  => mem_array(2)(84),
      output(3)  => mem_array(3)(84),
      output(4)  => mem_array(4)(84),
      output(5)  => mem_array(5)(84),
      output(6)  => mem_array(6)(84),
      output(7)  => mem_array(7)(84),
      output(8)  => mem_array(8)(84),
      output(9)  => mem_array(9)(84),
      output(10) => mem_array(10)(84),
      output(11) => mem_array(11)(84),
      output(12) => mem_array(12)(84),
      output(13) => mem_array(13)(84),
      output(14) => mem_array(14)(84),
      output(15) => mem_array(15)(84),
      output(16) => mem_array(16)(84),
      output(17) => mem_array(17)(84),
      output(18) => mem_array(18)(84),
      output(19) => mem_array(19)(84),
      output(20) => mem_array(20)(84),
      output(21) => mem_array(21)(84),
      output(22) => mem_array(22)(84),
      output(23) => mem_array(23)(84),
      output(24) => mem_array(24)(84),
      output(25) => mem_array(25)(84),
      output(26) => mem_array(26)(84),
      output(27) => mem_array(27)(84),
      output(28) => mem_array(28)(84),
      output(29) => mem_array(29)(84),
      output(30) => mem_array(30)(84),
      output(31) => mem_array(31)(84),
      output(32) => mem_array(32)(84),
      output(33) => mem_array(33)(84),
      output(34) => mem_array(34)(84),
      output(35) => mem_array(35)(84)
      );
  rom85 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001000000001001101000001101010010")
    port map (
      enable_o   => mem_enable_lines(85),
      output(0)  => mem_array(0)(85),
      output(1)  => mem_array(1)(85),
      output(2)  => mem_array(2)(85),
      output(3)  => mem_array(3)(85),
      output(4)  => mem_array(4)(85),
      output(5)  => mem_array(5)(85),
      output(6)  => mem_array(6)(85),
      output(7)  => mem_array(7)(85),
      output(8)  => mem_array(8)(85),
      output(9)  => mem_array(9)(85),
      output(10) => mem_array(10)(85),
      output(11) => mem_array(11)(85),
      output(12) => mem_array(12)(85),
      output(13) => mem_array(13)(85),
      output(14) => mem_array(14)(85),
      output(15) => mem_array(15)(85),
      output(16) => mem_array(16)(85),
      output(17) => mem_array(17)(85),
      output(18) => mem_array(18)(85),
      output(19) => mem_array(19)(85),
      output(20) => mem_array(20)(85),
      output(21) => mem_array(21)(85),
      output(22) => mem_array(22)(85),
      output(23) => mem_array(23)(85),
      output(24) => mem_array(24)(85),
      output(25) => mem_array(25)(85),
      output(26) => mem_array(26)(85),
      output(27) => mem_array(27)(85),
      output(28) => mem_array(28)(85),
      output(29) => mem_array(29)(85),
      output(30) => mem_array(30)(85),
      output(31) => mem_array(31)(85),
      output(32) => mem_array(32)(85),
      output(33) => mem_array(33)(85),
      output(34) => mem_array(34)(85),
      output(35) => mem_array(35)(85)
      );
  rom86 : entity work.rom
    generic map (
      bits  => 36,
      value => "000010000111000000100111000000110101")
    port map (
      enable_o   => mem_enable_lines(86),
      output(0)  => mem_array(0)(86),
      output(1)  => mem_array(1)(86),
      output(2)  => mem_array(2)(86),
      output(3)  => mem_array(3)(86),
      output(4)  => mem_array(4)(86),
      output(5)  => mem_array(5)(86),
      output(6)  => mem_array(6)(86),
      output(7)  => mem_array(7)(86),
      output(8)  => mem_array(8)(86),
      output(9)  => mem_array(9)(86),
      output(10) => mem_array(10)(86),
      output(11) => mem_array(11)(86),
      output(12) => mem_array(12)(86),
      output(13) => mem_array(13)(86),
      output(14) => mem_array(14)(86),
      output(15) => mem_array(15)(86),
      output(16) => mem_array(16)(86),
      output(17) => mem_array(17)(86),
      output(18) => mem_array(18)(86),
      output(19) => mem_array(19)(86),
      output(20) => mem_array(20)(86),
      output(21) => mem_array(21)(86),
      output(22) => mem_array(22)(86),
      output(23) => mem_array(23)(86),
      output(24) => mem_array(24)(86),
      output(25) => mem_array(25)(86),
      output(26) => mem_array(26)(86),
      output(27) => mem_array(27)(86),
      output(28) => mem_array(28)(86),
      output(29) => mem_array(29)(86),
      output(30) => mem_array(30)(86),
      output(31) => mem_array(31)(86),
      output(32) => mem_array(32)(86),
      output(33) => mem_array(33)(86),
      output(34) => mem_array(34)(86),
      output(35) => mem_array(35)(86)
      );
  rom87 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000100001000100000010011110001001")
    port map (
      enable_o   => mem_enable_lines(87),
      output(0)  => mem_array(0)(87),
      output(1)  => mem_array(1)(87),
      output(2)  => mem_array(2)(87),
      output(3)  => mem_array(3)(87),
      output(4)  => mem_array(4)(87),
      output(5)  => mem_array(5)(87),
      output(6)  => mem_array(6)(87),
      output(7)  => mem_array(7)(87),
      output(8)  => mem_array(8)(87),
      output(9)  => mem_array(9)(87),
      output(10) => mem_array(10)(87),
      output(11) => mem_array(11)(87),
      output(12) => mem_array(12)(87),
      output(13) => mem_array(13)(87),
      output(14) => mem_array(14)(87),
      output(15) => mem_array(15)(87),
      output(16) => mem_array(16)(87),
      output(17) => mem_array(17)(87),
      output(18) => mem_array(18)(87),
      output(19) => mem_array(19)(87),
      output(20) => mem_array(20)(87),
      output(21) => mem_array(21)(87),
      output(22) => mem_array(22)(87),
      output(23) => mem_array(23)(87),
      output(24) => mem_array(24)(87),
      output(25) => mem_array(25)(87),
      output(26) => mem_array(26)(87),
      output(27) => mem_array(27)(87),
      output(28) => mem_array(28)(87),
      output(29) => mem_array(29)(87),
      output(30) => mem_array(30)(87),
      output(31) => mem_array(31)(87),
      output(32) => mem_array(32)(87),
      output(33) => mem_array(33)(87),
      output(34) => mem_array(34)(87),
      output(35) => mem_array(35)(87)
      );
  rom88 : entity work.rom
    generic map (
      bits  => 36,
      value => "010010000000000000110000001010000000")
    port map (
      enable_o   => mem_enable_lines(88),
      output(0)  => mem_array(0)(88),
      output(1)  => mem_array(1)(88),
      output(2)  => mem_array(2)(88),
      output(3)  => mem_array(3)(88),
      output(4)  => mem_array(4)(88),
      output(5)  => mem_array(5)(88),
      output(6)  => mem_array(6)(88),
      output(7)  => mem_array(7)(88),
      output(8)  => mem_array(8)(88),
      output(9)  => mem_array(9)(88),
      output(10) => mem_array(10)(88),
      output(11) => mem_array(11)(88),
      output(12) => mem_array(12)(88),
      output(13) => mem_array(13)(88),
      output(14) => mem_array(14)(88),
      output(15) => mem_array(15)(88),
      output(16) => mem_array(16)(88),
      output(17) => mem_array(17)(88),
      output(18) => mem_array(18)(88),
      output(19) => mem_array(19)(88),
      output(20) => mem_array(20)(88),
      output(21) => mem_array(21)(88),
      output(22) => mem_array(22)(88),
      output(23) => mem_array(23)(88),
      output(24) => mem_array(24)(88),
      output(25) => mem_array(25)(88),
      output(26) => mem_array(26)(88),
      output(27) => mem_array(27)(88),
      output(28) => mem_array(28)(88),
      output(29) => mem_array(29)(88),
      output(30) => mem_array(30)(88),
      output(31) => mem_array(31)(88),
      output(32) => mem_array(32)(88),
      output(33) => mem_array(33)(88),
      output(34) => mem_array(34)(88),
      output(35) => mem_array(35)(88)
      );
  rom89 : entity work.rom
    generic map (
      bits  => 36,
      value => "000111001000000000000011000000101000")
    port map (
      enable_o   => mem_enable_lines(89),
      output(0)  => mem_array(0)(89),
      output(1)  => mem_array(1)(89),
      output(2)  => mem_array(2)(89),
      output(3)  => mem_array(3)(89),
      output(4)  => mem_array(4)(89),
      output(5)  => mem_array(5)(89),
      output(6)  => mem_array(6)(89),
      output(7)  => mem_array(7)(89),
      output(8)  => mem_array(8)(89),
      output(9)  => mem_array(9)(89),
      output(10) => mem_array(10)(89),
      output(11) => mem_array(11)(89),
      output(12) => mem_array(12)(89),
      output(13) => mem_array(13)(89),
      output(14) => mem_array(14)(89),
      output(15) => mem_array(15)(89),
      output(16) => mem_array(16)(89),
      output(17) => mem_array(17)(89),
      output(18) => mem_array(18)(89),
      output(19) => mem_array(19)(89),
      output(20) => mem_array(20)(89),
      output(21) => mem_array(21)(89),
      output(22) => mem_array(22)(89),
      output(23) => mem_array(23)(89),
      output(24) => mem_array(24)(89),
      output(25) => mem_array(25)(89),
      output(26) => mem_array(26)(89),
      output(27) => mem_array(27)(89),
      output(28) => mem_array(28)(89),
      output(29) => mem_array(29)(89),
      output(30) => mem_array(30)(89),
      output(31) => mem_array(31)(89),
      output(32) => mem_array(32)(89),
      output(33) => mem_array(33)(89),
      output(34) => mem_array(34)(89),
      output(35) => mem_array(35)(89)
      );
  rom90 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000111101000000010100010000000010")
    port map (
      enable_o   => mem_enable_lines(90),
      output(0)  => mem_array(0)(90),
      output(1)  => mem_array(1)(90),
      output(2)  => mem_array(2)(90),
      output(3)  => mem_array(3)(90),
      output(4)  => mem_array(4)(90),
      output(5)  => mem_array(5)(90),
      output(6)  => mem_array(6)(90),
      output(7)  => mem_array(7)(90),
      output(8)  => mem_array(8)(90),
      output(9)  => mem_array(9)(90),
      output(10) => mem_array(10)(90),
      output(11) => mem_array(11)(90),
      output(12) => mem_array(12)(90),
      output(13) => mem_array(13)(90),
      output(14) => mem_array(14)(90),
      output(15) => mem_array(15)(90),
      output(16) => mem_array(16)(90),
      output(17) => mem_array(17)(90),
      output(18) => mem_array(18)(90),
      output(19) => mem_array(19)(90),
      output(20) => mem_array(20)(90),
      output(21) => mem_array(21)(90),
      output(22) => mem_array(22)(90),
      output(23) => mem_array(23)(90),
      output(24) => mem_array(24)(90),
      output(25) => mem_array(25)(90),
      output(26) => mem_array(26)(90),
      output(27) => mem_array(27)(90),
      output(28) => mem_array(28)(90),
      output(29) => mem_array(29)(90),
      output(30) => mem_array(30)(90),
      output(31) => mem_array(31)(90),
      output(32) => mem_array(32)(90),
      output(33) => mem_array(33)(90),
      output(34) => mem_array(34)(90),
      output(35) => mem_array(35)(90)
      );
  rom91 : entity work.rom
    generic map (
      bits  => 36,
      value => "100100000001010000000100100000000000")
    port map (
      enable_o   => mem_enable_lines(91),
      output(0)  => mem_array(0)(91),
      output(1)  => mem_array(1)(91),
      output(2)  => mem_array(2)(91),
      output(3)  => mem_array(3)(91),
      output(4)  => mem_array(4)(91),
      output(5)  => mem_array(5)(91),
      output(6)  => mem_array(6)(91),
      output(7)  => mem_array(7)(91),
      output(8)  => mem_array(8)(91),
      output(9)  => mem_array(9)(91),
      output(10) => mem_array(10)(91),
      output(11) => mem_array(11)(91),
      output(12) => mem_array(12)(91),
      output(13) => mem_array(13)(91),
      output(14) => mem_array(14)(91),
      output(15) => mem_array(15)(91),
      output(16) => mem_array(16)(91),
      output(17) => mem_array(17)(91),
      output(18) => mem_array(18)(91),
      output(19) => mem_array(19)(91),
      output(20) => mem_array(20)(91),
      output(21) => mem_array(21)(91),
      output(22) => mem_array(22)(91),
      output(23) => mem_array(23)(91),
      output(24) => mem_array(24)(91),
      output(25) => mem_array(25)(91),
      output(26) => mem_array(26)(91),
      output(27) => mem_array(27)(91),
      output(28) => mem_array(28)(91),
      output(29) => mem_array(29)(91),
      output(30) => mem_array(30)(91),
      output(31) => mem_array(31)(91),
      output(32) => mem_array(32)(91),
      output(33) => mem_array(33)(91),
      output(34) => mem_array(34)(91),
      output(35) => mem_array(35)(91)
      );
  rom92 : entity work.rom
    generic map (
      bits  => 36,
      value => "001010011000000101000000000101001000")
    port map (
      enable_o   => mem_enable_lines(92),
      output(0)  => mem_array(0)(92),
      output(1)  => mem_array(1)(92),
      output(2)  => mem_array(2)(92),
      output(3)  => mem_array(3)(92),
      output(4)  => mem_array(4)(92),
      output(5)  => mem_array(5)(92),
      output(6)  => mem_array(6)(92),
      output(7)  => mem_array(7)(92),
      output(8)  => mem_array(8)(92),
      output(9)  => mem_array(9)(92),
      output(10) => mem_array(10)(92),
      output(11) => mem_array(11)(92),
      output(12) => mem_array(12)(92),
      output(13) => mem_array(13)(92),
      output(14) => mem_array(14)(92),
      output(15) => mem_array(15)(92),
      output(16) => mem_array(16)(92),
      output(17) => mem_array(17)(92),
      output(18) => mem_array(18)(92),
      output(19) => mem_array(19)(92),
      output(20) => mem_array(20)(92),
      output(21) => mem_array(21)(92),
      output(22) => mem_array(22)(92),
      output(23) => mem_array(23)(92),
      output(24) => mem_array(24)(92),
      output(25) => mem_array(25)(92),
      output(26) => mem_array(26)(92),
      output(27) => mem_array(27)(92),
      output(28) => mem_array(28)(92),
      output(29) => mem_array(29)(92),
      output(30) => mem_array(30)(92),
      output(31) => mem_array(31)(92),
      output(32) => mem_array(32)(92),
      output(33) => mem_array(33)(92),
      output(34) => mem_array(34)(92),
      output(35) => mem_array(35)(92)
      );
  rom93 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000101010000000110101000001001000")
    port map (
      enable_o   => mem_enable_lines(93),
      output(0)  => mem_array(0)(93),
      output(1)  => mem_array(1)(93),
      output(2)  => mem_array(2)(93),
      output(3)  => mem_array(3)(93),
      output(4)  => mem_array(4)(93),
      output(5)  => mem_array(5)(93),
      output(6)  => mem_array(6)(93),
      output(7)  => mem_array(7)(93),
      output(8)  => mem_array(8)(93),
      output(9)  => mem_array(9)(93),
      output(10) => mem_array(10)(93),
      output(11) => mem_array(11)(93),
      output(12) => mem_array(12)(93),
      output(13) => mem_array(13)(93),
      output(14) => mem_array(14)(93),
      output(15) => mem_array(15)(93),
      output(16) => mem_array(16)(93),
      output(17) => mem_array(17)(93),
      output(18) => mem_array(18)(93),
      output(19) => mem_array(19)(93),
      output(20) => mem_array(20)(93),
      output(21) => mem_array(21)(93),
      output(22) => mem_array(22)(93),
      output(23) => mem_array(23)(93),
      output(24) => mem_array(24)(93),
      output(25) => mem_array(25)(93),
      output(26) => mem_array(26)(93),
      output(27) => mem_array(27)(93),
      output(28) => mem_array(28)(93),
      output(29) => mem_array(29)(93),
      output(30) => mem_array(30)(93),
      output(31) => mem_array(31)(93),
      output(32) => mem_array(32)(93),
      output(33) => mem_array(33)(93),
      output(34) => mem_array(34)(93),
      output(35) => mem_array(35)(93)
      );
  rom94 : entity work.rom
    generic map (
      bits  => 36,
      value => "010000000010101010000001010000000001")
    port map (
      enable_o   => mem_enable_lines(94),
      output(0)  => mem_array(0)(94),
      output(1)  => mem_array(1)(94),
      output(2)  => mem_array(2)(94),
      output(3)  => mem_array(3)(94),
      output(4)  => mem_array(4)(94),
      output(5)  => mem_array(5)(94),
      output(6)  => mem_array(6)(94),
      output(7)  => mem_array(7)(94),
      output(8)  => mem_array(8)(94),
      output(9)  => mem_array(9)(94),
      output(10) => mem_array(10)(94),
      output(11) => mem_array(11)(94),
      output(12) => mem_array(12)(94),
      output(13) => mem_array(13)(94),
      output(14) => mem_array(14)(94),
      output(15) => mem_array(15)(94),
      output(16) => mem_array(16)(94),
      output(17) => mem_array(17)(94),
      output(18) => mem_array(18)(94),
      output(19) => mem_array(19)(94),
      output(20) => mem_array(20)(94),
      output(21) => mem_array(21)(94),
      output(22) => mem_array(22)(94),
      output(23) => mem_array(23)(94),
      output(24) => mem_array(24)(94),
      output(25) => mem_array(25)(94),
      output(26) => mem_array(26)(94),
      output(27) => mem_array(27)(94),
      output(28) => mem_array(28)(94),
      output(29) => mem_array(29)(94),
      output(30) => mem_array(30)(94),
      output(31) => mem_array(31)(94),
      output(32) => mem_array(32)(94),
      output(33) => mem_array(33)(94),
      output(34) => mem_array(34)(94),
      output(35) => mem_array(35)(94)
      );
  rom95 : entity work.rom
    generic map (
      bits  => 36,
      value => "010001010000001010110000001101010000")
    port map (
      enable_o   => mem_enable_lines(95),
      output(0)  => mem_array(0)(95),
      output(1)  => mem_array(1)(95),
      output(2)  => mem_array(2)(95),
      output(3)  => mem_array(3)(95),
      output(4)  => mem_array(4)(95),
      output(5)  => mem_array(5)(95),
      output(6)  => mem_array(6)(95),
      output(7)  => mem_array(7)(95),
      output(8)  => mem_array(8)(95),
      output(9)  => mem_array(9)(95),
      output(10) => mem_array(10)(95),
      output(11) => mem_array(11)(95),
      output(12) => mem_array(12)(95),
      output(13) => mem_array(13)(95),
      output(14) => mem_array(14)(95),
      output(15) => mem_array(15)(95),
      output(16) => mem_array(16)(95),
      output(17) => mem_array(17)(95),
      output(18) => mem_array(18)(95),
      output(19) => mem_array(19)(95),
      output(20) => mem_array(20)(95),
      output(21) => mem_array(21)(95),
      output(22) => mem_array(22)(95),
      output(23) => mem_array(23)(95),
      output(24) => mem_array(24)(95),
      output(25) => mem_array(25)(95),
      output(26) => mem_array(26)(95),
      output(27) => mem_array(27)(95),
      output(28) => mem_array(28)(95),
      output(29) => mem_array(29)(95),
      output(30) => mem_array(30)(95),
      output(31) => mem_array(31)(95),
      output(32) => mem_array(32)(95),
      output(33) => mem_array(33)(95),
      output(34) => mem_array(34)(95),
      output(35) => mem_array(35)(95)
      );
  rom96 : entity work.rom
    generic map (
      bits  => 36,
      value => "001000010001000000000001000000010100")
    port map (
      enable_o   => mem_enable_lines(96),
      output(0)  => mem_array(0)(96),
      output(1)  => mem_array(1)(96),
      output(2)  => mem_array(2)(96),
      output(3)  => mem_array(3)(96),
      output(4)  => mem_array(4)(96),
      output(5)  => mem_array(5)(96),
      output(6)  => mem_array(6)(96),
      output(7)  => mem_array(7)(96),
      output(8)  => mem_array(8)(96),
      output(9)  => mem_array(9)(96),
      output(10) => mem_array(10)(96),
      output(11) => mem_array(11)(96),
      output(12) => mem_array(12)(96),
      output(13) => mem_array(13)(96),
      output(14) => mem_array(14)(96),
      output(15) => mem_array(15)(96),
      output(16) => mem_array(16)(96),
      output(17) => mem_array(17)(96),
      output(18) => mem_array(18)(96),
      output(19) => mem_array(19)(96),
      output(20) => mem_array(20)(96),
      output(21) => mem_array(21)(96),
      output(22) => mem_array(22)(96),
      output(23) => mem_array(23)(96),
      output(24) => mem_array(24)(96),
      output(25) => mem_array(25)(96),
      output(26) => mem_array(26)(96),
      output(27) => mem_array(27)(96),
      output(28) => mem_array(28)(96),
      output(29) => mem_array(29)(96),
      output(30) => mem_array(30)(96),
      output(31) => mem_array(31)(96),
      output(32) => mem_array(32)(96),
      output(33) => mem_array(33)(96),
      output(34) => mem_array(34)(96),
      output(35) => mem_array(35)(96)
      );
  rom97 : entity work.rom
    generic map (
      bits  => 36,
      value => "000010000000011100000000011000000011")
    port map (
      enable_o   => mem_enable_lines(97),
      output(0)  => mem_array(0)(97),
      output(1)  => mem_array(1)(97),
      output(2)  => mem_array(2)(97),
      output(3)  => mem_array(3)(97),
      output(4)  => mem_array(4)(97),
      output(5)  => mem_array(5)(97),
      output(6)  => mem_array(6)(97),
      output(7)  => mem_array(7)(97),
      output(8)  => mem_array(8)(97),
      output(9)  => mem_array(9)(97),
      output(10) => mem_array(10)(97),
      output(11) => mem_array(11)(97),
      output(12) => mem_array(12)(97),
      output(13) => mem_array(13)(97),
      output(14) => mem_array(14)(97),
      output(15) => mem_array(15)(97),
      output(16) => mem_array(16)(97),
      output(17) => mem_array(17)(97),
      output(18) => mem_array(18)(97),
      output(19) => mem_array(19)(97),
      output(20) => mem_array(20)(97),
      output(21) => mem_array(21)(97),
      output(22) => mem_array(22)(97),
      output(23) => mem_array(23)(97),
      output(24) => mem_array(24)(97),
      output(25) => mem_array(25)(97),
      output(26) => mem_array(26)(97),
      output(27) => mem_array(27)(97),
      output(28) => mem_array(28)(97),
      output(29) => mem_array(29)(97),
      output(30) => mem_array(30)(97),
      output(31) => mem_array(31)(97),
      output(32) => mem_array(32)(97),
      output(33) => mem_array(33)(97),
      output(34) => mem_array(34)(97),
      output(35) => mem_array(35)(97)
      );
  rom98 : entity work.rom
    generic map (
      bits  => 36,
      value => "011000000100101001000000001011010000")
    port map (
      enable_o   => mem_enable_lines(98),
      output(0)  => mem_array(0)(98),
      output(1)  => mem_array(1)(98),
      output(2)  => mem_array(2)(98),
      output(3)  => mem_array(3)(98),
      output(4)  => mem_array(4)(98),
      output(5)  => mem_array(5)(98),
      output(6)  => mem_array(6)(98),
      output(7)  => mem_array(7)(98),
      output(8)  => mem_array(8)(98),
      output(9)  => mem_array(9)(98),
      output(10) => mem_array(10)(98),
      output(11) => mem_array(11)(98),
      output(12) => mem_array(12)(98),
      output(13) => mem_array(13)(98),
      output(14) => mem_array(14)(98),
      output(15) => mem_array(15)(98),
      output(16) => mem_array(16)(98),
      output(17) => mem_array(17)(98),
      output(18) => mem_array(18)(98),
      output(19) => mem_array(19)(98),
      output(20) => mem_array(20)(98),
      output(21) => mem_array(21)(98),
      output(22) => mem_array(22)(98),
      output(23) => mem_array(23)(98),
      output(24) => mem_array(24)(98),
      output(25) => mem_array(25)(98),
      output(26) => mem_array(26)(98),
      output(27) => mem_array(27)(98),
      output(28) => mem_array(28)(98),
      output(29) => mem_array(29)(98),
      output(30) => mem_array(30)(98),
      output(31) => mem_array(31)(98),
      output(32) => mem_array(32)(98),
      output(33) => mem_array(33)(98),
      output(34) => mem_array(34)(98),
      output(35) => mem_array(35)(98)
      );
  rom99 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000101")
    port map (
      enable_o   => mem_enable_lines(99),
      output(0)  => mem_array(0)(99),
      output(1)  => mem_array(1)(99),
      output(2)  => mem_array(2)(99),
      output(3)  => mem_array(3)(99),
      output(4)  => mem_array(4)(99),
      output(5)  => mem_array(5)(99),
      output(6)  => mem_array(6)(99),
      output(7)  => mem_array(7)(99),
      output(8)  => mem_array(8)(99),
      output(9)  => mem_array(9)(99),
      output(10) => mem_array(10)(99),
      output(11) => mem_array(11)(99),
      output(12) => mem_array(12)(99),
      output(13) => mem_array(13)(99),
      output(14) => mem_array(14)(99),
      output(15) => mem_array(15)(99),
      output(16) => mem_array(16)(99),
      output(17) => mem_array(17)(99),
      output(18) => mem_array(18)(99),
      output(19) => mem_array(19)(99),
      output(20) => mem_array(20)(99),
      output(21) => mem_array(21)(99),
      output(22) => mem_array(22)(99),
      output(23) => mem_array(23)(99),
      output(24) => mem_array(24)(99),
      output(25) => mem_array(25)(99),
      output(26) => mem_array(26)(99),
      output(27) => mem_array(27)(99),
      output(28) => mem_array(28)(99),
      output(29) => mem_array(29)(99),
      output(30) => mem_array(30)(99),
      output(31) => mem_array(31)(99),
      output(32) => mem_array(32)(99),
      output(33) => mem_array(33)(99),
      output(34) => mem_array(34)(99),
      output(35) => mem_array(35)(99)
      );
  rom100 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000110101000001001000010000000010")
    port map (
      enable_o   => mem_enable_lines(100),
      output(0)  => mem_array(0)(100),
      output(1)  => mem_array(1)(100),
      output(2)  => mem_array(2)(100),
      output(3)  => mem_array(3)(100),
      output(4)  => mem_array(4)(100),
      output(5)  => mem_array(5)(100),
      output(6)  => mem_array(6)(100),
      output(7)  => mem_array(7)(100),
      output(8)  => mem_array(8)(100),
      output(9)  => mem_array(9)(100),
      output(10) => mem_array(10)(100),
      output(11) => mem_array(11)(100),
      output(12) => mem_array(12)(100),
      output(13) => mem_array(13)(100),
      output(14) => mem_array(14)(100),
      output(15) => mem_array(15)(100),
      output(16) => mem_array(16)(100),
      output(17) => mem_array(17)(100),
      output(18) => mem_array(18)(100),
      output(19) => mem_array(19)(100),
      output(20) => mem_array(20)(100),
      output(21) => mem_array(21)(100),
      output(22) => mem_array(22)(100),
      output(23) => mem_array(23)(100),
      output(24) => mem_array(24)(100),
      output(25) => mem_array(25)(100),
      output(26) => mem_array(26)(100),
      output(27) => mem_array(27)(100),
      output(28) => mem_array(28)(100),
      output(29) => mem_array(29)(100),
      output(30) => mem_array(30)(100),
      output(31) => mem_array(31)(100),
      output(32) => mem_array(32)(100),
      output(33) => mem_array(33)(100),
      output(34) => mem_array(34)(100),
      output(35) => mem_array(35)(100)
      );
  rom101 : entity work.rom
    generic map (
      bits  => 36,
      value => "110110000001010000001000101000000000")
    port map (
      enable_o   => mem_enable_lines(101),
      output(0)  => mem_array(0)(101),
      output(1)  => mem_array(1)(101),
      output(2)  => mem_array(2)(101),
      output(3)  => mem_array(3)(101),
      output(4)  => mem_array(4)(101),
      output(5)  => mem_array(5)(101),
      output(6)  => mem_array(6)(101),
      output(7)  => mem_array(7)(101),
      output(8)  => mem_array(8)(101),
      output(9)  => mem_array(9)(101),
      output(10) => mem_array(10)(101),
      output(11) => mem_array(11)(101),
      output(12) => mem_array(12)(101),
      output(13) => mem_array(13)(101),
      output(14) => mem_array(14)(101),
      output(15) => mem_array(15)(101),
      output(16) => mem_array(16)(101),
      output(17) => mem_array(17)(101),
      output(18) => mem_array(18)(101),
      output(19) => mem_array(19)(101),
      output(20) => mem_array(20)(101),
      output(21) => mem_array(21)(101),
      output(22) => mem_array(22)(101),
      output(23) => mem_array(23)(101),
      output(24) => mem_array(24)(101),
      output(25) => mem_array(25)(101),
      output(26) => mem_array(26)(101),
      output(27) => mem_array(27)(101),
      output(28) => mem_array(28)(101),
      output(29) => mem_array(29)(101),
      output(30) => mem_array(30)(101),
      output(31) => mem_array(31)(101),
      output(32) => mem_array(32)(101),
      output(33) => mem_array(33)(101),
      output(34) => mem_array(34)(101),
      output(35) => mem_array(35)(101)
      );
  rom102 : entity work.rom
    generic map (
      bits  => 36,
      value => "001011100000001101010000000010000101")
    port map (
      enable_o   => mem_enable_lines(102),
      output(0)  => mem_array(0)(102),
      output(1)  => mem_array(1)(102),
      output(2)  => mem_array(2)(102),
      output(3)  => mem_array(3)(102),
      output(4)  => mem_array(4)(102),
      output(5)  => mem_array(5)(102),
      output(6)  => mem_array(6)(102),
      output(7)  => mem_array(7)(102),
      output(8)  => mem_array(8)(102),
      output(9)  => mem_array(9)(102),
      output(10) => mem_array(10)(102),
      output(11) => mem_array(11)(102),
      output(12) => mem_array(12)(102),
      output(13) => mem_array(13)(102),
      output(14) => mem_array(14)(102),
      output(15) => mem_array(15)(102),
      output(16) => mem_array(16)(102),
      output(17) => mem_array(17)(102),
      output(18) => mem_array(18)(102),
      output(19) => mem_array(19)(102),
      output(20) => mem_array(20)(102),
      output(21) => mem_array(21)(102),
      output(22) => mem_array(22)(102),
      output(23) => mem_array(23)(102),
      output(24) => mem_array(24)(102),
      output(25) => mem_array(25)(102),
      output(26) => mem_array(26)(102),
      output(27) => mem_array(27)(102),
      output(28) => mem_array(28)(102),
      output(29) => mem_array(29)(102),
      output(30) => mem_array(30)(102),
      output(31) => mem_array(31)(102),
      output(32) => mem_array(32)(102),
      output(33) => mem_array(33)(102),
      output(34) => mem_array(34)(102),
      output(35) => mem_array(35)(102)
      );
  rom103 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000101110100000010100000000100011")
    port map (
      enable_o   => mem_enable_lines(103),
      output(0)  => mem_array(0)(103),
      output(1)  => mem_array(1)(103),
      output(2)  => mem_array(2)(103),
      output(3)  => mem_array(3)(103),
      output(4)  => mem_array(4)(103),
      output(5)  => mem_array(5)(103),
      output(6)  => mem_array(6)(103),
      output(7)  => mem_array(7)(103),
      output(8)  => mem_array(8)(103),
      output(9)  => mem_array(9)(103),
      output(10) => mem_array(10)(103),
      output(11) => mem_array(11)(103),
      output(12) => mem_array(12)(103),
      output(13) => mem_array(13)(103),
      output(14) => mem_array(14)(103),
      output(15) => mem_array(15)(103),
      output(16) => mem_array(16)(103),
      output(17) => mem_array(17)(103),
      output(18) => mem_array(18)(103),
      output(19) => mem_array(19)(103),
      output(20) => mem_array(20)(103),
      output(21) => mem_array(21)(103),
      output(22) => mem_array(22)(103),
      output(23) => mem_array(23)(103),
      output(24) => mem_array(24)(103),
      output(25) => mem_array(25)(103),
      output(26) => mem_array(26)(103),
      output(27) => mem_array(27)(103),
      output(28) => mem_array(28)(103),
      output(29) => mem_array(29)(103),
      output(30) => mem_array(30)(103),
      output(31) => mem_array(31)(103),
      output(32) => mem_array(32)(103),
      output(33) => mem_array(33)(103),
      output(34) => mem_array(34)(103),
      output(35) => mem_array(35)(103)
      );
  rom104 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000010111100000001010000000000")
    port map (
      enable_o   => mem_enable_lines(104),
      output(0)  => mem_array(0)(104),
      output(1)  => mem_array(1)(104),
      output(2)  => mem_array(2)(104),
      output(3)  => mem_array(3)(104),
      output(4)  => mem_array(4)(104),
      output(5)  => mem_array(5)(104),
      output(6)  => mem_array(6)(104),
      output(7)  => mem_array(7)(104),
      output(8)  => mem_array(8)(104),
      output(9)  => mem_array(9)(104),
      output(10) => mem_array(10)(104),
      output(11) => mem_array(11)(104),
      output(12) => mem_array(12)(104),
      output(13) => mem_array(13)(104),
      output(14) => mem_array(14)(104),
      output(15) => mem_array(15)(104),
      output(16) => mem_array(16)(104),
      output(17) => mem_array(17)(104),
      output(18) => mem_array(18)(104),
      output(19) => mem_array(19)(104),
      output(20) => mem_array(20)(104),
      output(21) => mem_array(21)(104),
      output(22) => mem_array(22)(104),
      output(23) => mem_array(23)(104),
      output(24) => mem_array(24)(104),
      output(25) => mem_array(25)(104),
      output(26) => mem_array(26)(104),
      output(27) => mem_array(27)(104),
      output(28) => mem_array(28)(104),
      output(29) => mem_array(29)(104),
      output(30) => mem_array(30)(104),
      output(31) => mem_array(31)(104),
      output(32) => mem_array(32)(104),
      output(33) => mem_array(33)(104),
      output(34) => mem_array(34)(104),
      output(35) => mem_array(35)(104)
      );
  rom105 : entity work.rom
    generic map (
      bits  => 36,
      value => "100001000000001100001000000101000000")
    port map (
      enable_o   => mem_enable_lines(105),
      output(0)  => mem_array(0)(105),
      output(1)  => mem_array(1)(105),
      output(2)  => mem_array(2)(105),
      output(3)  => mem_array(3)(105),
      output(4)  => mem_array(4)(105),
      output(5)  => mem_array(5)(105),
      output(6)  => mem_array(6)(105),
      output(7)  => mem_array(7)(105),
      output(8)  => mem_array(8)(105),
      output(9)  => mem_array(9)(105),
      output(10) => mem_array(10)(105),
      output(11) => mem_array(11)(105),
      output(12) => mem_array(12)(105),
      output(13) => mem_array(13)(105),
      output(14) => mem_array(14)(105),
      output(15) => mem_array(15)(105),
      output(16) => mem_array(16)(105),
      output(17) => mem_array(17)(105),
      output(18) => mem_array(18)(105),
      output(19) => mem_array(19)(105),
      output(20) => mem_array(20)(105),
      output(21) => mem_array(21)(105),
      output(22) => mem_array(22)(105),
      output(23) => mem_array(23)(105),
      output(24) => mem_array(24)(105),
      output(25) => mem_array(25)(105),
      output(26) => mem_array(26)(105),
      output(27) => mem_array(27)(105),
      output(28) => mem_array(28)(105),
      output(29) => mem_array(29)(105),
      output(30) => mem_array(30)(105),
      output(31) => mem_array(31)(105),
      output(32) => mem_array(32)(105),
      output(33) => mem_array(33)(105),
      output(34) => mem_array(34)(105),
      output(35) => mem_array(35)(105)
      );
  rom106 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000000000000000000111000000110110")
    port map (
      enable_o   => mem_enable_lines(106),
      output(0)  => mem_array(0)(106),
      output(1)  => mem_array(1)(106),
      output(2)  => mem_array(2)(106),
      output(3)  => mem_array(3)(106),
      output(4)  => mem_array(4)(106),
      output(5)  => mem_array(5)(106),
      output(6)  => mem_array(6)(106),
      output(7)  => mem_array(7)(106),
      output(8)  => mem_array(8)(106),
      output(9)  => mem_array(9)(106),
      output(10) => mem_array(10)(106),
      output(11) => mem_array(11)(106),
      output(12) => mem_array(12)(106),
      output(13) => mem_array(13)(106),
      output(14) => mem_array(14)(106),
      output(15) => mem_array(15)(106),
      output(16) => mem_array(16)(106),
      output(17) => mem_array(17)(106),
      output(18) => mem_array(18)(106),
      output(19) => mem_array(19)(106),
      output(20) => mem_array(20)(106),
      output(21) => mem_array(21)(106),
      output(22) => mem_array(22)(106),
      output(23) => mem_array(23)(106),
      output(24) => mem_array(24)(106),
      output(25) => mem_array(25)(106),
      output(26) => mem_array(26)(106),
      output(27) => mem_array(27)(106),
      output(28) => mem_array(28)(106),
      output(29) => mem_array(29)(106),
      output(30) => mem_array(30)(106),
      output(31) => mem_array(31)(106),
      output(32) => mem_array(32)(106),
      output(33) => mem_array(33)(106),
      output(34) => mem_array(34)(106),
      output(35) => mem_array(35)(106)
      );
  rom107 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001010010000000000000110000011")
    port map (
      enable_o   => mem_enable_lines(107),
      output(0)  => mem_array(0)(107),
      output(1)  => mem_array(1)(107),
      output(2)  => mem_array(2)(107),
      output(3)  => mem_array(3)(107),
      output(4)  => mem_array(4)(107),
      output(5)  => mem_array(5)(107),
      output(6)  => mem_array(6)(107),
      output(7)  => mem_array(7)(107),
      output(8)  => mem_array(8)(107),
      output(9)  => mem_array(9)(107),
      output(10) => mem_array(10)(107),
      output(11) => mem_array(11)(107),
      output(12) => mem_array(12)(107),
      output(13) => mem_array(13)(107),
      output(14) => mem_array(14)(107),
      output(15) => mem_array(15)(107),
      output(16) => mem_array(16)(107),
      output(17) => mem_array(17)(107),
      output(18) => mem_array(18)(107),
      output(19) => mem_array(19)(107),
      output(20) => mem_array(20)(107),
      output(21) => mem_array(21)(107),
      output(22) => mem_array(22)(107),
      output(23) => mem_array(23)(107),
      output(24) => mem_array(24)(107),
      output(25) => mem_array(25)(107),
      output(26) => mem_array(26)(107),
      output(27) => mem_array(27)(107),
      output(28) => mem_array(28)(107),
      output(29) => mem_array(29)(107),
      output(30) => mem_array(30)(107),
      output(31) => mem_array(31)(107),
      output(32) => mem_array(32)(107),
      output(33) => mem_array(33)(107),
      output(34) => mem_array(34)(107),
      output(35) => mem_array(35)(107)
      );
  rom108 : entity work.rom
    generic map (
      bits  => 36,
      value => "011000000100101001000000000000010000")
    port map (
      enable_o   => mem_enable_lines(108),
      output(0)  => mem_array(0)(108),
      output(1)  => mem_array(1)(108),
      output(2)  => mem_array(2)(108),
      output(3)  => mem_array(3)(108),
      output(4)  => mem_array(4)(108),
      output(5)  => mem_array(5)(108),
      output(6)  => mem_array(6)(108),
      output(7)  => mem_array(7)(108),
      output(8)  => mem_array(8)(108),
      output(9)  => mem_array(9)(108),
      output(10) => mem_array(10)(108),
      output(11) => mem_array(11)(108),
      output(12) => mem_array(12)(108),
      output(13) => mem_array(13)(108),
      output(14) => mem_array(14)(108),
      output(15) => mem_array(15)(108),
      output(16) => mem_array(16)(108),
      output(17) => mem_array(17)(108),
      output(18) => mem_array(18)(108),
      output(19) => mem_array(19)(108),
      output(20) => mem_array(20)(108),
      output(21) => mem_array(21)(108),
      output(22) => mem_array(22)(108),
      output(23) => mem_array(23)(108),
      output(24) => mem_array(24)(108),
      output(25) => mem_array(25)(108),
      output(26) => mem_array(26)(108),
      output(27) => mem_array(27)(108),
      output(28) => mem_array(28)(108),
      output(29) => mem_array(29)(108),
      output(30) => mem_array(30)(108),
      output(31) => mem_array(31)(108),
      output(32) => mem_array(32)(108),
      output(33) => mem_array(33)(108),
      output(34) => mem_array(34)(108),
      output(35) => mem_array(35)(108)
      );
  rom109 : entity work.rom
    generic map (
      bits  => 36,
      value => "000101000000000101000111000000110001")
    port map (
      enable_o   => mem_enable_lines(109),
      output(0)  => mem_array(0)(109),
      output(1)  => mem_array(1)(109),
      output(2)  => mem_array(2)(109),
      output(3)  => mem_array(3)(109),
      output(4)  => mem_array(4)(109),
      output(5)  => mem_array(5)(109),
      output(6)  => mem_array(6)(109),
      output(7)  => mem_array(7)(109),
      output(8)  => mem_array(8)(109),
      output(9)  => mem_array(9)(109),
      output(10) => mem_array(10)(109),
      output(11) => mem_array(11)(109),
      output(12) => mem_array(12)(109),
      output(13) => mem_array(13)(109),
      output(14) => mem_array(14)(109),
      output(15) => mem_array(15)(109),
      output(16) => mem_array(16)(109),
      output(17) => mem_array(17)(109),
      output(18) => mem_array(18)(109),
      output(19) => mem_array(19)(109),
      output(20) => mem_array(20)(109),
      output(21) => mem_array(21)(109),
      output(22) => mem_array(22)(109),
      output(23) => mem_array(23)(109),
      output(24) => mem_array(24)(109),
      output(25) => mem_array(25)(109),
      output(26) => mem_array(26)(109),
      output(27) => mem_array(27)(109),
      output(28) => mem_array(28)(109),
      output(29) => mem_array(29)(109),
      output(30) => mem_array(30)(109),
      output(31) => mem_array(31)(109),
      output(32) => mem_array(32)(109),
      output(33) => mem_array(33)(109),
      output(34) => mem_array(34)(109),
      output(35) => mem_array(35)(109)
      );
  rom110 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000111100010000000000100000000011")
    port map (
      enable_o   => mem_enable_lines(110),
      output(0)  => mem_array(0)(110),
      output(1)  => mem_array(1)(110),
      output(2)  => mem_array(2)(110),
      output(3)  => mem_array(3)(110),
      output(4)  => mem_array(4)(110),
      output(5)  => mem_array(5)(110),
      output(6)  => mem_array(6)(110),
      output(7)  => mem_array(7)(110),
      output(8)  => mem_array(8)(110),
      output(9)  => mem_array(9)(110),
      output(10) => mem_array(10)(110),
      output(11) => mem_array(11)(110),
      output(12) => mem_array(12)(110),
      output(13) => mem_array(13)(110),
      output(14) => mem_array(14)(110),
      output(15) => mem_array(15)(110),
      output(16) => mem_array(16)(110),
      output(17) => mem_array(17)(110),
      output(18) => mem_array(18)(110),
      output(19) => mem_array(19)(110),
      output(20) => mem_array(20)(110),
      output(21) => mem_array(21)(110),
      output(22) => mem_array(22)(110),
      output(23) => mem_array(23)(110),
      output(24) => mem_array(24)(110),
      output(25) => mem_array(25)(110),
      output(26) => mem_array(26)(110),
      output(27) => mem_array(27)(110),
      output(28) => mem_array(28)(110),
      output(29) => mem_array(29)(110),
      output(30) => mem_array(30)(110),
      output(31) => mem_array(31)(110),
      output(32) => mem_array(32)(110),
      output(33) => mem_array(33)(110),
      output(34) => mem_array(34)(110),
      output(35) => mem_array(35)(110)
      );
  rom111 : entity work.rom
    generic map (
      bits  => 36,
      value => "001010000011110000000000100010000000")
    port map (
      enable_o   => mem_enable_lines(111),
      output(0)  => mem_array(0)(111),
      output(1)  => mem_array(1)(111),
      output(2)  => mem_array(2)(111),
      output(3)  => mem_array(3)(111),
      output(4)  => mem_array(4)(111),
      output(5)  => mem_array(5)(111),
      output(6)  => mem_array(6)(111),
      output(7)  => mem_array(7)(111),
      output(8)  => mem_array(8)(111),
      output(9)  => mem_array(9)(111),
      output(10) => mem_array(10)(111),
      output(11) => mem_array(11)(111),
      output(12) => mem_array(12)(111),
      output(13) => mem_array(13)(111),
      output(14) => mem_array(14)(111),
      output(15) => mem_array(15)(111),
      output(16) => mem_array(16)(111),
      output(17) => mem_array(17)(111),
      output(18) => mem_array(18)(111),
      output(19) => mem_array(19)(111),
      output(20) => mem_array(20)(111),
      output(21) => mem_array(21)(111),
      output(22) => mem_array(22)(111),
      output(23) => mem_array(23)(111),
      output(24) => mem_array(24)(111),
      output(25) => mem_array(25)(111),
      output(26) => mem_array(26)(111),
      output(27) => mem_array(27)(111),
      output(28) => mem_array(28)(111),
      output(29) => mem_array(29)(111),
      output(30) => mem_array(30)(111),
      output(31) => mem_array(31)(111),
      output(32) => mem_array(32)(111),
      output(33) => mem_array(33)(111),
      output(34) => mem_array(34)(111),
      output(35) => mem_array(35)(111)
      );
  rom112 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000101000001101100000010010100100")
    port map (
      enable_o   => mem_enable_lines(112),
      output(0)  => mem_array(0)(112),
      output(1)  => mem_array(1)(112),
      output(2)  => mem_array(2)(112),
      output(3)  => mem_array(3)(112),
      output(4)  => mem_array(4)(112),
      output(5)  => mem_array(5)(112),
      output(6)  => mem_array(6)(112),
      output(7)  => mem_array(7)(112),
      output(8)  => mem_array(8)(112),
      output(9)  => mem_array(9)(112),
      output(10) => mem_array(10)(112),
      output(11) => mem_array(11)(112),
      output(12) => mem_array(12)(112),
      output(13) => mem_array(13)(112),
      output(14) => mem_array(14)(112),
      output(15) => mem_array(15)(112),
      output(16) => mem_array(16)(112),
      output(17) => mem_array(17)(112),
      output(18) => mem_array(18)(112),
      output(19) => mem_array(19)(112),
      output(20) => mem_array(20)(112),
      output(21) => mem_array(21)(112),
      output(22) => mem_array(22)(112),
      output(23) => mem_array(23)(112),
      output(24) => mem_array(24)(112),
      output(25) => mem_array(25)(112),
      output(26) => mem_array(26)(112),
      output(27) => mem_array(27)(112),
      output(28) => mem_array(28)(112),
      output(29) => mem_array(29)(112),
      output(30) => mem_array(30)(112),
      output(31) => mem_array(31)(112),
      output(32) => mem_array(32)(112),
      output(33) => mem_array(33)(112),
      output(34) => mem_array(34)(112),
      output(35) => mem_array(35)(112)
      );
  rom113 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000110011000000010001110000000000")
    port map (
      enable_o   => mem_enable_lines(113),
      output(0)  => mem_array(0)(113),
      output(1)  => mem_array(1)(113),
      output(2)  => mem_array(2)(113),
      output(3)  => mem_array(3)(113),
      output(4)  => mem_array(4)(113),
      output(5)  => mem_array(5)(113),
      output(6)  => mem_array(6)(113),
      output(7)  => mem_array(7)(113),
      output(8)  => mem_array(8)(113),
      output(9)  => mem_array(9)(113),
      output(10) => mem_array(10)(113),
      output(11) => mem_array(11)(113),
      output(12) => mem_array(12)(113),
      output(13) => mem_array(13)(113),
      output(14) => mem_array(14)(113),
      output(15) => mem_array(15)(113),
      output(16) => mem_array(16)(113),
      output(17) => mem_array(17)(113),
      output(18) => mem_array(18)(113),
      output(19) => mem_array(19)(113),
      output(20) => mem_array(20)(113),
      output(21) => mem_array(21)(113),
      output(22) => mem_array(22)(113),
      output(23) => mem_array(23)(113),
      output(24) => mem_array(24)(113),
      output(25) => mem_array(25)(113),
      output(26) => mem_array(26)(113),
      output(27) => mem_array(27)(113),
      output(28) => mem_array(28)(113),
      output(29) => mem_array(29)(113),
      output(30) => mem_array(30)(113),
      output(31) => mem_array(31)(113),
      output(32) => mem_array(32)(113),
      output(33) => mem_array(33)(113),
      output(34) => mem_array(34)(113),
      output(35) => mem_array(35)(113)
      );
  rom114 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000011001110000011110011000000")
    port map (
      enable_o   => mem_enable_lines(114),
      output(0)  => mem_array(0)(114),
      output(1)  => mem_array(1)(114),
      output(2)  => mem_array(2)(114),
      output(3)  => mem_array(3)(114),
      output(4)  => mem_array(4)(114),
      output(5)  => mem_array(5)(114),
      output(6)  => mem_array(6)(114),
      output(7)  => mem_array(7)(114),
      output(8)  => mem_array(8)(114),
      output(9)  => mem_array(9)(114),
      output(10) => mem_array(10)(114),
      output(11) => mem_array(11)(114),
      output(12) => mem_array(12)(114),
      output(13) => mem_array(13)(114),
      output(14) => mem_array(14)(114),
      output(15) => mem_array(15)(114),
      output(16) => mem_array(16)(114),
      output(17) => mem_array(17)(114),
      output(18) => mem_array(18)(114),
      output(19) => mem_array(19)(114),
      output(20) => mem_array(20)(114),
      output(21) => mem_array(21)(114),
      output(22) => mem_array(22)(114),
      output(23) => mem_array(23)(114),
      output(24) => mem_array(24)(114),
      output(25) => mem_array(25)(114),
      output(26) => mem_array(26)(114),
      output(27) => mem_array(27)(114),
      output(28) => mem_array(28)(114),
      output(29) => mem_array(29)(114),
      output(30) => mem_array(30)(114),
      output(31) => mem_array(31)(114),
      output(32) => mem_array(32)(114),
      output(33) => mem_array(33)(114),
      output(34) => mem_array(34)(114),
      output(35) => mem_array(35)(114)
      );
  rom115 : entity work.rom
    generic map (
      bits  => 36,
      value => "000010000000001101000000001111001100")
    port map (
      enable_o   => mem_enable_lines(115),
      output(0)  => mem_array(0)(115),
      output(1)  => mem_array(1)(115),
      output(2)  => mem_array(2)(115),
      output(3)  => mem_array(3)(115),
      output(4)  => mem_array(4)(115),
      output(5)  => mem_array(5)(115),
      output(6)  => mem_array(6)(115),
      output(7)  => mem_array(7)(115),
      output(8)  => mem_array(8)(115),
      output(9)  => mem_array(9)(115),
      output(10) => mem_array(10)(115),
      output(11) => mem_array(11)(115),
      output(12) => mem_array(12)(115),
      output(13) => mem_array(13)(115),
      output(14) => mem_array(14)(115),
      output(15) => mem_array(15)(115),
      output(16) => mem_array(16)(115),
      output(17) => mem_array(17)(115),
      output(18) => mem_array(18)(115),
      output(19) => mem_array(19)(115),
      output(20) => mem_array(20)(115),
      output(21) => mem_array(21)(115),
      output(22) => mem_array(22)(115),
      output(23) => mem_array(23)(115),
      output(24) => mem_array(24)(115),
      output(25) => mem_array(25)(115),
      output(26) => mem_array(26)(115),
      output(27) => mem_array(27)(115),
      output(28) => mem_array(28)(115),
      output(29) => mem_array(29)(115),
      output(30) => mem_array(30)(115),
      output(31) => mem_array(31)(115),
      output(32) => mem_array(32)(115),
      output(33) => mem_array(33)(115),
      output(34) => mem_array(34)(115),
      output(35) => mem_array(35)(115)
      );
  rom116 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001000000000110100100000111100")
    port map (
      enable_o   => mem_enable_lines(116),
      output(0)  => mem_array(0)(116),
      output(1)  => mem_array(1)(116),
      output(2)  => mem_array(2)(116),
      output(3)  => mem_array(3)(116),
      output(4)  => mem_array(4)(116),
      output(5)  => mem_array(5)(116),
      output(6)  => mem_array(6)(116),
      output(7)  => mem_array(7)(116),
      output(8)  => mem_array(8)(116),
      output(9)  => mem_array(9)(116),
      output(10) => mem_array(10)(116),
      output(11) => mem_array(11)(116),
      output(12) => mem_array(12)(116),
      output(13) => mem_array(13)(116),
      output(14) => mem_array(14)(116),
      output(15) => mem_array(15)(116),
      output(16) => mem_array(16)(116),
      output(17) => mem_array(17)(116),
      output(18) => mem_array(18)(116),
      output(19) => mem_array(19)(116),
      output(20) => mem_array(20)(116),
      output(21) => mem_array(21)(116),
      output(22) => mem_array(22)(116),
      output(23) => mem_array(23)(116),
      output(24) => mem_array(24)(116),
      output(25) => mem_array(25)(116),
      output(26) => mem_array(26)(116),
      output(27) => mem_array(27)(116),
      output(28) => mem_array(28)(116),
      output(29) => mem_array(29)(116),
      output(30) => mem_array(30)(116),
      output(31) => mem_array(31)(116),
      output(32) => mem_array(32)(116),
      output(33) => mem_array(33)(116),
      output(34) => mem_array(34)(116),
      output(35) => mem_array(35)(116)
      );
  rom117 : entity work.rom
    generic map (
      bits  => 36,
      value => "110000000000100000000011010100000011")
    port map (
      enable_o   => mem_enable_lines(117),
      output(0)  => mem_array(0)(117),
      output(1)  => mem_array(1)(117),
      output(2)  => mem_array(2)(117),
      output(3)  => mem_array(3)(117),
      output(4)  => mem_array(4)(117),
      output(5)  => mem_array(5)(117),
      output(6)  => mem_array(6)(117),
      output(7)  => mem_array(7)(117),
      output(8)  => mem_array(8)(117),
      output(9)  => mem_array(9)(117),
      output(10) => mem_array(10)(117),
      output(11) => mem_array(11)(117),
      output(12) => mem_array(12)(117),
      output(13) => mem_array(13)(117),
      output(14) => mem_array(14)(117),
      output(15) => mem_array(15)(117),
      output(16) => mem_array(16)(117),
      output(17) => mem_array(17)(117),
      output(18) => mem_array(18)(117),
      output(19) => mem_array(19)(117),
      output(20) => mem_array(20)(117),
      output(21) => mem_array(21)(117),
      output(22) => mem_array(22)(117),
      output(23) => mem_array(23)(117),
      output(24) => mem_array(24)(117),
      output(25) => mem_array(25)(117),
      output(26) => mem_array(26)(117),
      output(27) => mem_array(27)(117),
      output(28) => mem_array(28)(117),
      output(29) => mem_array(29)(117),
      output(30) => mem_array(30)(117),
      output(31) => mem_array(31)(117),
      output(32) => mem_array(32)(117),
      output(33) => mem_array(33)(117),
      output(34) => mem_array(34)(117),
      output(35) => mem_array(35)(117)
      );
  rom118 : entity work.rom
    generic map (
      bits  => 36,
      value => "110111000000000010000000001101011000")
    port map (
      enable_o   => mem_enable_lines(118),
      output(0)  => mem_array(0)(118),
      output(1)  => mem_array(1)(118),
      output(2)  => mem_array(2)(118),
      output(3)  => mem_array(3)(118),
      output(4)  => mem_array(4)(118),
      output(5)  => mem_array(5)(118),
      output(6)  => mem_array(6)(118),
      output(7)  => mem_array(7)(118),
      output(8)  => mem_array(8)(118),
      output(9)  => mem_array(9)(118),
      output(10) => mem_array(10)(118),
      output(11) => mem_array(11)(118),
      output(12) => mem_array(12)(118),
      output(13) => mem_array(13)(118),
      output(14) => mem_array(14)(118),
      output(15) => mem_array(15)(118),
      output(16) => mem_array(16)(118),
      output(17) => mem_array(17)(118),
      output(18) => mem_array(18)(118),
      output(19) => mem_array(19)(118),
      output(20) => mem_array(20)(118),
      output(21) => mem_array(21)(118),
      output(22) => mem_array(22)(118),
      output(23) => mem_array(23)(118),
      output(24) => mem_array(24)(118),
      output(25) => mem_array(25)(118),
      output(26) => mem_array(26)(118),
      output(27) => mem_array(27)(118),
      output(28) => mem_array(28)(118),
      output(29) => mem_array(29)(118),
      output(30) => mem_array(30)(118),
      output(31) => mem_array(31)(118),
      output(32) => mem_array(32)(118),
      output(33) => mem_array(33)(118),
      output(34) => mem_array(34)(118),
      output(35) => mem_array(35)(118)
      );
  rom119 : entity work.rom
    generic map (
      bits  => 36,
      value => "001111001100000000001000000000110110")
    port map (
      enable_o   => mem_enable_lines(119),
      output(0)  => mem_array(0)(119),
      output(1)  => mem_array(1)(119),
      output(2)  => mem_array(2)(119),
      output(3)  => mem_array(3)(119),
      output(4)  => mem_array(4)(119),
      output(5)  => mem_array(5)(119),
      output(6)  => mem_array(6)(119),
      output(7)  => mem_array(7)(119),
      output(8)  => mem_array(8)(119),
      output(9)  => mem_array(9)(119),
      output(10) => mem_array(10)(119),
      output(11) => mem_array(11)(119),
      output(12) => mem_array(12)(119),
      output(13) => mem_array(13)(119),
      output(14) => mem_array(14)(119),
      output(15) => mem_array(15)(119),
      output(16) => mem_array(16)(119),
      output(17) => mem_array(17)(119),
      output(18) => mem_array(18)(119),
      output(19) => mem_array(19)(119),
      output(20) => mem_array(20)(119),
      output(21) => mem_array(21)(119),
      output(22) => mem_array(22)(119),
      output(23) => mem_array(23)(119),
      output(24) => mem_array(24)(119),
      output(25) => mem_array(25)(119),
      output(26) => mem_array(26)(119),
      output(27) => mem_array(27)(119),
      output(28) => mem_array(28)(119),
      output(29) => mem_array(29)(119),
      output(30) => mem_array(30)(119),
      output(31) => mem_array(31)(119),
      output(32) => mem_array(32)(119),
      output(33) => mem_array(33)(119),
      output(34) => mem_array(34)(119),
      output(35) => mem_array(35)(119)
      );
  rom120 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000111101000000010100100000000011")
    port map (
      enable_o   => mem_enable_lines(120),
      output(0)  => mem_array(0)(120),
      output(1)  => mem_array(1)(120),
      output(2)  => mem_array(2)(120),
      output(3)  => mem_array(3)(120),
      output(4)  => mem_array(4)(120),
      output(5)  => mem_array(5)(120),
      output(6)  => mem_array(6)(120),
      output(7)  => mem_array(7)(120),
      output(8)  => mem_array(8)(120),
      output(9)  => mem_array(9)(120),
      output(10) => mem_array(10)(120),
      output(11) => mem_array(11)(120),
      output(12) => mem_array(12)(120),
      output(13) => mem_array(13)(120),
      output(14) => mem_array(14)(120),
      output(15) => mem_array(15)(120),
      output(16) => mem_array(16)(120),
      output(17) => mem_array(17)(120),
      output(18) => mem_array(18)(120),
      output(19) => mem_array(19)(120),
      output(20) => mem_array(20)(120),
      output(21) => mem_array(21)(120),
      output(22) => mem_array(22)(120),
      output(23) => mem_array(23)(120),
      output(24) => mem_array(24)(120),
      output(25) => mem_array(25)(120),
      output(26) => mem_array(26)(120),
      output(27) => mem_array(27)(120),
      output(28) => mem_array(28)(120),
      output(29) => mem_array(29)(120),
      output(30) => mem_array(30)(120),
      output(31) => mem_array(31)(120),
      output(32) => mem_array(32)(120),
      output(33) => mem_array(33)(120),
      output(34) => mem_array(34)(120),
      output(35) => mem_array(35)(120)
      );
  rom121 : entity work.rom
    generic map (
      bits  => 36,
      value => "011010000001000111000000000000000000")
    port map (
      enable_o   => mem_enable_lines(121),
      output(0)  => mem_array(0)(121),
      output(1)  => mem_array(1)(121),
      output(2)  => mem_array(2)(121),
      output(3)  => mem_array(3)(121),
      output(4)  => mem_array(4)(121),
      output(5)  => mem_array(5)(121),
      output(6)  => mem_array(6)(121),
      output(7)  => mem_array(7)(121),
      output(8)  => mem_array(8)(121),
      output(9)  => mem_array(9)(121),
      output(10) => mem_array(10)(121),
      output(11) => mem_array(11)(121),
      output(12) => mem_array(12)(121),
      output(13) => mem_array(13)(121),
      output(14) => mem_array(14)(121),
      output(15) => mem_array(15)(121),
      output(16) => mem_array(16)(121),
      output(17) => mem_array(17)(121),
      output(18) => mem_array(18)(121),
      output(19) => mem_array(19)(121),
      output(20) => mem_array(20)(121),
      output(21) => mem_array(21)(121),
      output(22) => mem_array(22)(121),
      output(23) => mem_array(23)(121),
      output(24) => mem_array(24)(121),
      output(25) => mem_array(25)(121),
      output(26) => mem_array(26)(121),
      output(27) => mem_array(27)(121),
      output(28) => mem_array(28)(121),
      output(29) => mem_array(29)(121),
      output(30) => mem_array(30)(121),
      output(31) => mem_array(31)(121),
      output(32) => mem_array(32)(121),
      output(33) => mem_array(33)(121),
      output(34) => mem_array(34)(121),
      output(35) => mem_array(35)(121)
      );
  rom122 : entity work.rom
    generic map (
      bits  => 36,
      value => "001101110000001111001100000000001000")
    port map (
      enable_o   => mem_enable_lines(122),
      output(0)  => mem_array(0)(122),
      output(1)  => mem_array(1)(122),
      output(2)  => mem_array(2)(122),
      output(3)  => mem_array(3)(122),
      output(4)  => mem_array(4)(122),
      output(5)  => mem_array(5)(122),
      output(6)  => mem_array(6)(122),
      output(7)  => mem_array(7)(122),
      output(8)  => mem_array(8)(122),
      output(9)  => mem_array(9)(122),
      output(10) => mem_array(10)(122),
      output(11) => mem_array(11)(122),
      output(12) => mem_array(12)(122),
      output(13) => mem_array(13)(122),
      output(14) => mem_array(14)(122),
      output(15) => mem_array(15)(122),
      output(16) => mem_array(16)(122),
      output(17) => mem_array(17)(122),
      output(18) => mem_array(18)(122),
      output(19) => mem_array(19)(122),
      output(20) => mem_array(20)(122),
      output(21) => mem_array(21)(122),
      output(22) => mem_array(22)(122),
      output(23) => mem_array(23)(122),
      output(24) => mem_array(24)(122),
      output(25) => mem_array(25)(122),
      output(26) => mem_array(26)(122),
      output(27) => mem_array(27)(122),
      output(28) => mem_array(28)(122),
      output(29) => mem_array(29)(122),
      output(30) => mem_array(30)(122),
      output(31) => mem_array(31)(122),
      output(32) => mem_array(32)(122),
      output(33) => mem_array(33)(122),
      output(34) => mem_array(34)(122),
      output(35) => mem_array(35)(122)
      );
  rom123 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000110111100000111101110000000000")
    port map (
      enable_o   => mem_enable_lines(123),
      output(0)  => mem_array(0)(123),
      output(1)  => mem_array(1)(123),
      output(2)  => mem_array(2)(123),
      output(3)  => mem_array(3)(123),
      output(4)  => mem_array(4)(123),
      output(5)  => mem_array(5)(123),
      output(6)  => mem_array(6)(123),
      output(7)  => mem_array(7)(123),
      output(8)  => mem_array(8)(123),
      output(9)  => mem_array(9)(123),
      output(10) => mem_array(10)(123),
      output(11) => mem_array(11)(123),
      output(12) => mem_array(12)(123),
      output(13) => mem_array(13)(123),
      output(14) => mem_array(14)(123),
      output(15) => mem_array(15)(123),
      output(16) => mem_array(16)(123),
      output(17) => mem_array(17)(123),
      output(18) => mem_array(18)(123),
      output(19) => mem_array(19)(123),
      output(20) => mem_array(20)(123),
      output(21) => mem_array(21)(123),
      output(22) => mem_array(22)(123),
      output(23) => mem_array(23)(123),
      output(24) => mem_array(24)(123),
      output(25) => mem_array(25)(123),
      output(26) => mem_array(26)(123),
      output(27) => mem_array(27)(123),
      output(28) => mem_array(28)(123),
      output(29) => mem_array(29)(123),
      output(30) => mem_array(30)(123),
      output(31) => mem_array(31)(123),
      output(32) => mem_array(32)(123),
      output(33) => mem_array(33)(123),
      output(34) => mem_array(34)(123),
      output(35) => mem_array(35)(123)
      );
  rom124 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000000011100000000011110011000000")
    port map (
      enable_o   => mem_enable_lines(124),
      output(0)  => mem_array(0)(124),
      output(1)  => mem_array(1)(124),
      output(2)  => mem_array(2)(124),
      output(3)  => mem_array(3)(124),
      output(4)  => mem_array(4)(124),
      output(5)  => mem_array(5)(124),
      output(6)  => mem_array(6)(124),
      output(7)  => mem_array(7)(124),
      output(8)  => mem_array(8)(124),
      output(9)  => mem_array(9)(124),
      output(10) => mem_array(10)(124),
      output(11) => mem_array(11)(124),
      output(12) => mem_array(12)(124),
      output(13) => mem_array(13)(124),
      output(14) => mem_array(14)(124),
      output(15) => mem_array(15)(124),
      output(16) => mem_array(16)(124),
      output(17) => mem_array(17)(124),
      output(18) => mem_array(18)(124),
      output(19) => mem_array(19)(124),
      output(20) => mem_array(20)(124),
      output(21) => mem_array(21)(124),
      output(22) => mem_array(22)(124),
      output(23) => mem_array(23)(124),
      output(24) => mem_array(24)(124),
      output(25) => mem_array(25)(124),
      output(26) => mem_array(26)(124),
      output(27) => mem_array(27)(124),
      output(28) => mem_array(28)(124),
      output(29) => mem_array(29)(124),
      output(30) => mem_array(30)(124),
      output(31) => mem_array(31)(124),
      output(32) => mem_array(32)(124),
      output(33) => mem_array(33)(124),
      output(34) => mem_array(34)(124),
      output(35) => mem_array(35)(124)
      );
  rom125 : entity work.rom
    generic map (
      bits  => 36,
      value => "000010000000001110001000001111001100")
    port map (
      enable_o   => mem_enable_lines(125),
      output(0)  => mem_array(0)(125),
      output(1)  => mem_array(1)(125),
      output(2)  => mem_array(2)(125),
      output(3)  => mem_array(3)(125),
      output(4)  => mem_array(4)(125),
      output(5)  => mem_array(5)(125),
      output(6)  => mem_array(6)(125),
      output(7)  => mem_array(7)(125),
      output(8)  => mem_array(8)(125),
      output(9)  => mem_array(9)(125),
      output(10) => mem_array(10)(125),
      output(11) => mem_array(11)(125),
      output(12) => mem_array(12)(125),
      output(13) => mem_array(13)(125),
      output(14) => mem_array(14)(125),
      output(15) => mem_array(15)(125),
      output(16) => mem_array(16)(125),
      output(17) => mem_array(17)(125),
      output(18) => mem_array(18)(125),
      output(19) => mem_array(19)(125),
      output(20) => mem_array(20)(125),
      output(21) => mem_array(21)(125),
      output(22) => mem_array(22)(125),
      output(23) => mem_array(23)(125),
      output(24) => mem_array(24)(125),
      output(25) => mem_array(25)(125),
      output(26) => mem_array(26)(125),
      output(27) => mem_array(27)(125),
      output(28) => mem_array(28)(125),
      output(29) => mem_array(29)(125),
      output(30) => mem_array(30)(125),
      output(31) => mem_array(31)(125),
      output(32) => mem_array(32)(125),
      output(33) => mem_array(33)(125),
      output(34) => mem_array(34)(125),
      output(35) => mem_array(35)(125)
      );
  rom126 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001000000000111001000000111101")
    port map (
      enable_o   => mem_enable_lines(126),
      output(0)  => mem_array(0)(126),
      output(1)  => mem_array(1)(126),
      output(2)  => mem_array(2)(126),
      output(3)  => mem_array(3)(126),
      output(4)  => mem_array(4)(126),
      output(5)  => mem_array(5)(126),
      output(6)  => mem_array(6)(126),
      output(7)  => mem_array(7)(126),
      output(8)  => mem_array(8)(126),
      output(9)  => mem_array(9)(126),
      output(10) => mem_array(10)(126),
      output(11) => mem_array(11)(126),
      output(12) => mem_array(12)(126),
      output(13) => mem_array(13)(126),
      output(14) => mem_array(14)(126),
      output(15) => mem_array(15)(126),
      output(16) => mem_array(16)(126),
      output(17) => mem_array(17)(126),
      output(18) => mem_array(18)(126),
      output(19) => mem_array(19)(126),
      output(20) => mem_array(20)(126),
      output(21) => mem_array(21)(126),
      output(22) => mem_array(22)(126),
      output(23) => mem_array(23)(126),
      output(24) => mem_array(24)(126),
      output(25) => mem_array(25)(126),
      output(26) => mem_array(26)(126),
      output(27) => mem_array(27)(126),
      output(28) => mem_array(28)(126),
      output(29) => mem_array(29)(126),
      output(30) => mem_array(30)(126),
      output(31) => mem_array(31)(126),
      output(32) => mem_array(32)(126),
      output(33) => mem_array(33)(126),
      output(34) => mem_array(34)(126),
      output(35) => mem_array(35)(126)
      );
  rom127 : entity work.rom
    generic map (
      bits  => 36,
      value => "110000000000100000000011100110000011")
    port map (
      enable_o   => mem_enable_lines(127),
      output(0)  => mem_array(0)(127),
      output(1)  => mem_array(1)(127),
      output(2)  => mem_array(2)(127),
      output(3)  => mem_array(3)(127),
      output(4)  => mem_array(4)(127),
      output(5)  => mem_array(5)(127),
      output(6)  => mem_array(6)(127),
      output(7)  => mem_array(7)(127),
      output(8)  => mem_array(8)(127),
      output(9)  => mem_array(9)(127),
      output(10) => mem_array(10)(127),
      output(11) => mem_array(11)(127),
      output(12) => mem_array(12)(127),
      output(13) => mem_array(13)(127),
      output(14) => mem_array(14)(127),
      output(15) => mem_array(15)(127),
      output(16) => mem_array(16)(127),
      output(17) => mem_array(17)(127),
      output(18) => mem_array(18)(127),
      output(19) => mem_array(19)(127),
      output(20) => mem_array(20)(127),
      output(21) => mem_array(21)(127),
      output(22) => mem_array(22)(127),
      output(23) => mem_array(23)(127),
      output(24) => mem_array(24)(127),
      output(25) => mem_array(25)(127),
      output(26) => mem_array(26)(127),
      output(27) => mem_array(27)(127),
      output(28) => mem_array(28)(127),
      output(29) => mem_array(29)(127),
      output(30) => mem_array(30)(127),
      output(31) => mem_array(31)(127),
      output(32) => mem_array(32)(127),
      output(33) => mem_array(33)(127),
      output(34) => mem_array(34)(127),
      output(35) => mem_array(35)(127)
      );
  rom128 : entity work.rom
    generic map (
      bits  => 36,
      value => "110000000001010010000000001110100000")
    port map (
      enable_o   => mem_enable_lines(128),
      output(0)  => mem_array(0)(128),
      output(1)  => mem_array(1)(128),
      output(2)  => mem_array(2)(128),
      output(3)  => mem_array(3)(128),
      output(4)  => mem_array(4)(128),
      output(5)  => mem_array(5)(128),
      output(6)  => mem_array(6)(128),
      output(7)  => mem_array(7)(128),
      output(8)  => mem_array(8)(128),
      output(9)  => mem_array(9)(128),
      output(10) => mem_array(10)(128),
      output(11) => mem_array(11)(128),
      output(12) => mem_array(12)(128),
      output(13) => mem_array(13)(128),
      output(14) => mem_array(14)(128),
      output(15) => mem_array(15)(128),
      output(16) => mem_array(16)(128),
      output(17) => mem_array(17)(128),
      output(18) => mem_array(18)(128),
      output(19) => mem_array(19)(128),
      output(20) => mem_array(20)(128),
      output(21) => mem_array(21)(128),
      output(22) => mem_array(22)(128),
      output(23) => mem_array(23)(128),
      output(24) => mem_array(24)(128),
      output(25) => mem_array(25)(128),
      output(26) => mem_array(26)(128),
      output(27) => mem_array(27)(128),
      output(28) => mem_array(28)(128),
      output(29) => mem_array(29)(128),
      output(30) => mem_array(30)(128),
      output(31) => mem_array(31)(128),
      output(32) => mem_array(32)(128),
      output(33) => mem_array(33)(128),
      output(34) => mem_array(34)(128),
      output(35) => mem_array(35)(128)
      );
  rom129 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000111010")
    port map (
      enable_o   => mem_enable_lines(129),
      output(0)  => mem_array(0)(129),
      output(1)  => mem_array(1)(129),
      output(2)  => mem_array(2)(129),
      output(3)  => mem_array(3)(129),
      output(4)  => mem_array(4)(129),
      output(5)  => mem_array(5)(129),
      output(6)  => mem_array(6)(129),
      output(7)  => mem_array(7)(129),
      output(8)  => mem_array(8)(129),
      output(9)  => mem_array(9)(129),
      output(10) => mem_array(10)(129),
      output(11) => mem_array(11)(129),
      output(12) => mem_array(12)(129),
      output(13) => mem_array(13)(129),
      output(14) => mem_array(14)(129),
      output(15) => mem_array(15)(129),
      output(16) => mem_array(16)(129),
      output(17) => mem_array(17)(129),
      output(18) => mem_array(18)(129),
      output(19) => mem_array(19)(129),
      output(20) => mem_array(20)(129),
      output(21) => mem_array(21)(129),
      output(22) => mem_array(22)(129),
      output(23) => mem_array(23)(129),
      output(24) => mem_array(24)(129),
      output(25) => mem_array(25)(129),
      output(26) => mem_array(26)(129),
      output(27) => mem_array(27)(129),
      output(28) => mem_array(28)(129),
      output(29) => mem_array(29)(129),
      output(30) => mem_array(30)(129),
      output(31) => mem_array(31)(129),
      output(32) => mem_array(32)(129),
      output(33) => mem_array(33)(129),
      output(34) => mem_array(34)(129),
      output(35) => mem_array(35)(129)
      );
  rom130 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000111100000000010100100000000011")
    port map (
      enable_o   => mem_enable_lines(130),
      output(0)  => mem_array(0)(130),
      output(1)  => mem_array(1)(130),
      output(2)  => mem_array(2)(130),
      output(3)  => mem_array(3)(130),
      output(4)  => mem_array(4)(130),
      output(5)  => mem_array(5)(130),
      output(6)  => mem_array(6)(130),
      output(7)  => mem_array(7)(130),
      output(8)  => mem_array(8)(130),
      output(9)  => mem_array(9)(130),
      output(10) => mem_array(10)(130),
      output(11) => mem_array(11)(130),
      output(12) => mem_array(12)(130),
      output(13) => mem_array(13)(130),
      output(14) => mem_array(14)(130),
      output(15) => mem_array(15)(130),
      output(16) => mem_array(16)(130),
      output(17) => mem_array(17)(130),
      output(18) => mem_array(18)(130),
      output(19) => mem_array(19)(130),
      output(20) => mem_array(20)(130),
      output(21) => mem_array(21)(130),
      output(22) => mem_array(22)(130),
      output(23) => mem_array(23)(130),
      output(24) => mem_array(24)(130),
      output(25) => mem_array(25)(130),
      output(26) => mem_array(26)(130),
      output(27) => mem_array(27)(130),
      output(28) => mem_array(28)(130),
      output(29) => mem_array(29)(130),
      output(30) => mem_array(30)(130),
      output(31) => mem_array(31)(130),
      output(32) => mem_array(32)(130),
      output(33) => mem_array(33)(130),
      output(34) => mem_array(34)(130),
      output(35) => mem_array(35)(130)
      );
  rom131 : entity work.rom
    generic map (
      bits  => 36,
      value => "101100000001000111000000000000000000")
    port map (
      enable_o   => mem_enable_lines(131),
      output(0)  => mem_array(0)(131),
      output(1)  => mem_array(1)(131),
      output(2)  => mem_array(2)(131),
      output(3)  => mem_array(3)(131),
      output(4)  => mem_array(4)(131),
      output(5)  => mem_array(5)(131),
      output(6)  => mem_array(6)(131),
      output(7)  => mem_array(7)(131),
      output(8)  => mem_array(8)(131),
      output(9)  => mem_array(9)(131),
      output(10) => mem_array(10)(131),
      output(11) => mem_array(11)(131),
      output(12) => mem_array(12)(131),
      output(13) => mem_array(13)(131),
      output(14) => mem_array(14)(131),
      output(15) => mem_array(15)(131),
      output(16) => mem_array(16)(131),
      output(17) => mem_array(17)(131),
      output(18) => mem_array(18)(131),
      output(19) => mem_array(19)(131),
      output(20) => mem_array(20)(131),
      output(21) => mem_array(21)(131),
      output(22) => mem_array(22)(131),
      output(23) => mem_array(23)(131),
      output(24) => mem_array(24)(131),
      output(25) => mem_array(25)(131),
      output(26) => mem_array(26)(131),
      output(27) => mem_array(27)(131),
      output(28) => mem_array(28)(131),
      output(29) => mem_array(29)(131),
      output(30) => mem_array(30)(131),
      output(31) => mem_array(31)(131),
      output(32) => mem_array(32)(131),
      output(33) => mem_array(33)(131),
      output(34) => mem_array(34)(131),
      output(35) => mem_array(35)(131)
      );
  rom132 : entity work.rom
    generic map (
      bits  => 36,
      value => "001110111000001111001100000000001000")
    port map (
      enable_o   => mem_enable_lines(132),
      output(0)  => mem_array(0)(132),
      output(1)  => mem_array(1)(132),
      output(2)  => mem_array(2)(132),
      output(3)  => mem_array(3)(132),
      output(4)  => mem_array(4)(132),
      output(5)  => mem_array(5)(132),
      output(6)  => mem_array(6)(132),
      output(7)  => mem_array(7)(132),
      output(8)  => mem_array(8)(132),
      output(9)  => mem_array(9)(132),
      output(10) => mem_array(10)(132),
      output(11) => mem_array(11)(132),
      output(12) => mem_array(12)(132),
      output(13) => mem_array(13)(132),
      output(14) => mem_array(14)(132),
      output(15) => mem_array(15)(132),
      output(16) => mem_array(16)(132),
      output(17) => mem_array(17)(132),
      output(18) => mem_array(18)(132),
      output(19) => mem_array(19)(132),
      output(20) => mem_array(20)(132),
      output(21) => mem_array(21)(132),
      output(22) => mem_array(22)(132),
      output(23) => mem_array(23)(132),
      output(24) => mem_array(24)(132),
      output(25) => mem_array(25)(132),
      output(26) => mem_array(26)(132),
      output(27) => mem_array(27)(132),
      output(28) => mem_array(28)(132),
      output(29) => mem_array(29)(132),
      output(30) => mem_array(30)(132),
      output(31) => mem_array(31)(132),
      output(32) => mem_array(32)(132),
      output(33) => mem_array(33)(132),
      output(34) => mem_array(34)(132),
      output(35) => mem_array(35)(132)
      );
  rom133 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000111100000000111100110000000000")
    port map (
      enable_o   => mem_enable_lines(133),
      output(0)  => mem_array(0)(133),
      output(1)  => mem_array(1)(133),
      output(2)  => mem_array(2)(133),
      output(3)  => mem_array(3)(133),
      output(4)  => mem_array(4)(133),
      output(5)  => mem_array(5)(133),
      output(6)  => mem_array(6)(133),
      output(7)  => mem_array(7)(133),
      output(8)  => mem_array(8)(133),
      output(9)  => mem_array(9)(133),
      output(10) => mem_array(10)(133),
      output(11) => mem_array(11)(133),
      output(12) => mem_array(12)(133),
      output(13) => mem_array(13)(133),
      output(14) => mem_array(14)(133),
      output(15) => mem_array(15)(133),
      output(16) => mem_array(16)(133),
      output(17) => mem_array(17)(133),
      output(18) => mem_array(18)(133),
      output(19) => mem_array(19)(133),
      output(20) => mem_array(20)(133),
      output(21) => mem_array(21)(133),
      output(22) => mem_array(22)(133),
      output(23) => mem_array(23)(133),
      output(24) => mem_array(24)(133),
      output(25) => mem_array(25)(133),
      output(26) => mem_array(26)(133),
      output(27) => mem_array(27)(133),
      output(28) => mem_array(28)(133),
      output(29) => mem_array(29)(133),
      output(30) => mem_array(30)(133),
      output(31) => mem_array(31)(133),
      output(32) => mem_array(32)(133),
      output(33) => mem_array(33)(133),
      output(34) => mem_array(34)(133),
      output(35) => mem_array(35)(133)
      );
  rom134 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000000011110010000011110111000000")
    port map (
      enable_o   => mem_enable_lines(134),
      output(0)  => mem_array(0)(134),
      output(1)  => mem_array(1)(134),
      output(2)  => mem_array(2)(134),
      output(3)  => mem_array(3)(134),
      output(4)  => mem_array(4)(134),
      output(5)  => mem_array(5)(134),
      output(6)  => mem_array(6)(134),
      output(7)  => mem_array(7)(134),
      output(8)  => mem_array(8)(134),
      output(9)  => mem_array(9)(134),
      output(10) => mem_array(10)(134),
      output(11) => mem_array(11)(134),
      output(12) => mem_array(12)(134),
      output(13) => mem_array(13)(134),
      output(14) => mem_array(14)(134),
      output(15) => mem_array(15)(134),
      output(16) => mem_array(16)(134),
      output(17) => mem_array(17)(134),
      output(18) => mem_array(18)(134),
      output(19) => mem_array(19)(134),
      output(20) => mem_array(20)(134),
      output(21) => mem_array(21)(134),
      output(22) => mem_array(22)(134),
      output(23) => mem_array(23)(134),
      output(24) => mem_array(24)(134),
      output(25) => mem_array(25)(134),
      output(26) => mem_array(26)(134),
      output(27) => mem_array(27)(134),
      output(28) => mem_array(28)(134),
      output(29) => mem_array(29)(134),
      output(30) => mem_array(30)(134),
      output(31) => mem_array(31)(134),
      output(32) => mem_array(32)(134),
      output(33) => mem_array(33)(134),
      output(34) => mem_array(34)(134),
      output(35) => mem_array(35)(134)
      );
  rom135 : entity work.rom
    generic map (
      bits  => 36,
      value => "000010000000001111010000001111011100")
    port map (
      enable_o   => mem_enable_lines(135),
      output(0)  => mem_array(0)(135),
      output(1)  => mem_array(1)(135),
      output(2)  => mem_array(2)(135),
      output(3)  => mem_array(3)(135),
      output(4)  => mem_array(4)(135),
      output(5)  => mem_array(5)(135),
      output(6)  => mem_array(6)(135),
      output(7)  => mem_array(7)(135),
      output(8)  => mem_array(8)(135),
      output(9)  => mem_array(9)(135),
      output(10) => mem_array(10)(135),
      output(11) => mem_array(11)(135),
      output(12) => mem_array(12)(135),
      output(13) => mem_array(13)(135),
      output(14) => mem_array(14)(135),
      output(15) => mem_array(15)(135),
      output(16) => mem_array(16)(135),
      output(17) => mem_array(17)(135),
      output(18) => mem_array(18)(135),
      output(19) => mem_array(19)(135),
      output(20) => mem_array(20)(135),
      output(21) => mem_array(21)(135),
      output(22) => mem_array(22)(135),
      output(23) => mem_array(23)(135),
      output(24) => mem_array(24)(135),
      output(25) => mem_array(25)(135),
      output(26) => mem_array(26)(135),
      output(27) => mem_array(27)(135),
      output(28) => mem_array(28)(135),
      output(29) => mem_array(29)(135),
      output(30) => mem_array(30)(135),
      output(31) => mem_array(31)(135),
      output(32) => mem_array(32)(135),
      output(33) => mem_array(33)(135),
      output(34) => mem_array(34)(135),
      output(35) => mem_array(35)(135)
      );
  rom136 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001000000000111101100000111101")
    port map (
      enable_o   => mem_enable_lines(136),
      output(0)  => mem_array(0)(136),
      output(1)  => mem_array(1)(136),
      output(2)  => mem_array(2)(136),
      output(3)  => mem_array(3)(136),
      output(4)  => mem_array(4)(136),
      output(5)  => mem_array(5)(136),
      output(6)  => mem_array(6)(136),
      output(7)  => mem_array(7)(136),
      output(8)  => mem_array(8)(136),
      output(9)  => mem_array(9)(136),
      output(10) => mem_array(10)(136),
      output(11) => mem_array(11)(136),
      output(12) => mem_array(12)(136),
      output(13) => mem_array(13)(136),
      output(14) => mem_array(14)(136),
      output(15) => mem_array(15)(136),
      output(16) => mem_array(16)(136),
      output(17) => mem_array(17)(136),
      output(18) => mem_array(18)(136),
      output(19) => mem_array(19)(136),
      output(20) => mem_array(20)(136),
      output(21) => mem_array(21)(136),
      output(22) => mem_array(22)(136),
      output(23) => mem_array(23)(136),
      output(24) => mem_array(24)(136),
      output(25) => mem_array(25)(136),
      output(26) => mem_array(26)(136),
      output(27) => mem_array(27)(136),
      output(28) => mem_array(28)(136),
      output(29) => mem_array(29)(136),
      output(30) => mem_array(30)(136),
      output(31) => mem_array(31)(136),
      output(32) => mem_array(32)(136),
      output(33) => mem_array(33)(136),
      output(34) => mem_array(34)(136),
      output(35) => mem_array(35)(136)
      );
  rom137 : entity work.rom
    generic map (
      bits  => 36,
      value => "110000000000100000000011111000000011")
    port map (
      enable_o   => mem_enable_lines(137),
      output(0)  => mem_array(0)(137),
      output(1)  => mem_array(1)(137),
      output(2)  => mem_array(2)(137),
      output(3)  => mem_array(3)(137),
      output(4)  => mem_array(4)(137),
      output(5)  => mem_array(5)(137),
      output(6)  => mem_array(6)(137),
      output(7)  => mem_array(7)(137),
      output(8)  => mem_array(8)(137),
      output(9)  => mem_array(9)(137),
      output(10) => mem_array(10)(137),
      output(11) => mem_array(11)(137),
      output(12) => mem_array(12)(137),
      output(13) => mem_array(13)(137),
      output(14) => mem_array(14)(137),
      output(15) => mem_array(15)(137),
      output(16) => mem_array(16)(137),
      output(17) => mem_array(17)(137),
      output(18) => mem_array(18)(137),
      output(19) => mem_array(19)(137),
      output(20) => mem_array(20)(137),
      output(21) => mem_array(21)(137),
      output(22) => mem_array(22)(137),
      output(23) => mem_array(23)(137),
      output(24) => mem_array(24)(137),
      output(25) => mem_array(25)(137),
      output(26) => mem_array(26)(137),
      output(27) => mem_array(27)(137),
      output(28) => mem_array(28)(137),
      output(29) => mem_array(29)(137),
      output(30) => mem_array(30)(137),
      output(31) => mem_array(31)(137),
      output(32) => mem_array(32)(137),
      output(33) => mem_array(33)(137),
      output(34) => mem_array(34)(137),
      output(35) => mem_array(35)(137)
      );
  rom138 : entity work.rom
    generic map (
      bits  => 36,
      value => "110100000001010010000000001111101000")
    port map (
      enable_o   => mem_enable_lines(138),
      output(0)  => mem_array(0)(138),
      output(1)  => mem_array(1)(138),
      output(2)  => mem_array(2)(138),
      output(3)  => mem_array(3)(138),
      output(4)  => mem_array(4)(138),
      output(5)  => mem_array(5)(138),
      output(6)  => mem_array(6)(138),
      output(7)  => mem_array(7)(138),
      output(8)  => mem_array(8)(138),
      output(9)  => mem_array(9)(138),
      output(10) => mem_array(10)(138),
      output(11) => mem_array(11)(138),
      output(12) => mem_array(12)(138),
      output(13) => mem_array(13)(138),
      output(14) => mem_array(14)(138),
      output(15) => mem_array(15)(138),
      output(16) => mem_array(16)(138),
      output(17) => mem_array(17)(138),
      output(18) => mem_array(18)(138),
      output(19) => mem_array(19)(138),
      output(20) => mem_array(20)(138),
      output(21) => mem_array(21)(138),
      output(22) => mem_array(22)(138),
      output(23) => mem_array(23)(138),
      output(24) => mem_array(24)(138),
      output(25) => mem_array(25)(138),
      output(26) => mem_array(26)(138),
      output(27) => mem_array(27)(138),
      output(28) => mem_array(28)(138),
      output(29) => mem_array(29)(138),
      output(30) => mem_array(30)(138),
      output(31) => mem_array(31)(138),
      output(32) => mem_array(32)(138),
      output(33) => mem_array(33)(138),
      output(34) => mem_array(34)(138),
      output(35) => mem_array(35)(138)
      );
  rom139 : entity work.rom
    generic map (
      bits  => 36,
      value => "000100011100000000000000000000111111")
    port map (
      enable_o   => mem_enable_lines(139),
      output(0)  => mem_array(0)(139),
      output(1)  => mem_array(1)(139),
      output(2)  => mem_array(2)(139),
      output(3)  => mem_array(3)(139),
      output(4)  => mem_array(4)(139),
      output(5)  => mem_array(5)(139),
      output(6)  => mem_array(6)(139),
      output(7)  => mem_array(7)(139),
      output(8)  => mem_array(8)(139),
      output(9)  => mem_array(9)(139),
      output(10) => mem_array(10)(139),
      output(11) => mem_array(11)(139),
      output(12) => mem_array(12)(139),
      output(13) => mem_array(13)(139),
      output(14) => mem_array(14)(139),
      output(15) => mem_array(15)(139),
      output(16) => mem_array(16)(139),
      output(17) => mem_array(17)(139),
      output(18) => mem_array(18)(139),
      output(19) => mem_array(19)(139),
      output(20) => mem_array(20)(139),
      output(21) => mem_array(21)(139),
      output(22) => mem_array(22)(139),
      output(23) => mem_array(23)(139),
      output(24) => mem_array(24)(139),
      output(25) => mem_array(25)(139),
      output(26) => mem_array(26)(139),
      output(27) => mem_array(27)(139),
      output(28) => mem_array(28)(139),
      output(29) => mem_array(29)(139),
      output(30) => mem_array(30)(139),
      output(31) => mem_array(31)(139),
      output(32) => mem_array(32)(139),
      output(33) => mem_array(33)(139),
      output(34) => mem_array(34)(139),
      output(35) => mem_array(35)(139)
      );
  rom140 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000111100110000000000100000000000")
    port map (
      enable_o   => mem_enable_lines(140),
      output(0)  => mem_array(0)(140),
      output(1)  => mem_array(1)(140),
      output(2)  => mem_array(2)(140),
      output(3)  => mem_array(3)(140),
      output(4)  => mem_array(4)(140),
      output(5)  => mem_array(5)(140),
      output(6)  => mem_array(6)(140),
      output(7)  => mem_array(7)(140),
      output(8)  => mem_array(8)(140),
      output(9)  => mem_array(9)(140),
      output(10) => mem_array(10)(140),
      output(11) => mem_array(11)(140),
      output(12) => mem_array(12)(140),
      output(13) => mem_array(13)(140),
      output(14) => mem_array(14)(140),
      output(15) => mem_array(15)(140),
      output(16) => mem_array(16)(140),
      output(17) => mem_array(17)(140),
      output(18) => mem_array(18)(140),
      output(19) => mem_array(19)(140),
      output(20) => mem_array(20)(140),
      output(21) => mem_array(21)(140),
      output(22) => mem_array(22)(140),
      output(23) => mem_array(23)(140),
      output(24) => mem_array(24)(140),
      output(25) => mem_array(25)(140),
      output(26) => mem_array(26)(140),
      output(27) => mem_array(27)(140),
      output(28) => mem_array(28)(140),
      output(29) => mem_array(29)(140),
      output(30) => mem_array(30)(140),
      output(31) => mem_array(31)(140),
      output(32) => mem_array(32)(140),
      output(33) => mem_array(33)(140),
      output(34) => mem_array(34)(140),
      output(35) => mem_array(35)(140)
      );
  rom141 : entity work.rom
    generic map (
      bits  => 36,
      value => "001110000011011000000100101001000000")
    port map (
      enable_o   => mem_enable_lines(141),
      output(0)  => mem_array(0)(141),
      output(1)  => mem_array(1)(141),
      output(2)  => mem_array(2)(141),
      output(3)  => mem_array(3)(141),
      output(4)  => mem_array(4)(141),
      output(5)  => mem_array(5)(141),
      output(6)  => mem_array(6)(141),
      output(7)  => mem_array(7)(141),
      output(8)  => mem_array(8)(141),
      output(9)  => mem_array(9)(141),
      output(10) => mem_array(10)(141),
      output(11) => mem_array(11)(141),
      output(12) => mem_array(12)(141),
      output(13) => mem_array(13)(141),
      output(14) => mem_array(14)(141),
      output(15) => mem_array(15)(141),
      output(16) => mem_array(16)(141),
      output(17) => mem_array(17)(141),
      output(18) => mem_array(18)(141),
      output(19) => mem_array(19)(141),
      output(20) => mem_array(20)(141),
      output(21) => mem_array(21)(141),
      output(22) => mem_array(22)(141),
      output(23) => mem_array(23)(141),
      output(24) => mem_array(24)(141),
      output(25) => mem_array(25)(141),
      output(26) => mem_array(26)(141),
      output(27) => mem_array(27)(141),
      output(28) => mem_array(28)(141),
      output(29) => mem_array(29)(141),
      output(30) => mem_array(30)(141),
      output(31) => mem_array(31)(141),
      output(32) => mem_array(32)(141),
      output(33) => mem_array(33)(141),
      output(34) => mem_array(34)(141),
      output(35) => mem_array(35)(141)
      );
  rom142 : entity work.rom
    generic map (
      bits  => 36,
      value => "010000000000001111011100000000001000")
    port map (
      enable_o   => mem_enable_lines(142),
      output(0)  => mem_array(0)(142),
      output(1)  => mem_array(1)(142),
      output(2)  => mem_array(2)(142),
      output(3)  => mem_array(3)(142),
      output(4)  => mem_array(4)(142),
      output(5)  => mem_array(5)(142),
      output(6)  => mem_array(6)(142),
      output(7)  => mem_array(7)(142),
      output(8)  => mem_array(8)(142),
      output(9)  => mem_array(9)(142),
      output(10) => mem_array(10)(142),
      output(11) => mem_array(11)(142),
      output(12) => mem_array(12)(142),
      output(13) => mem_array(13)(142),
      output(14) => mem_array(14)(142),
      output(15) => mem_array(15)(142),
      output(16) => mem_array(16)(142),
      output(17) => mem_array(17)(142),
      output(18) => mem_array(18)(142),
      output(19) => mem_array(19)(142),
      output(20) => mem_array(20)(142),
      output(21) => mem_array(21)(142),
      output(22) => mem_array(22)(142),
      output(23) => mem_array(23)(142),
      output(24) => mem_array(24)(142),
      output(25) => mem_array(25)(142),
      output(26) => mem_array(26)(142),
      output(27) => mem_array(27)(142),
      output(28) => mem_array(28)(142),
      output(29) => mem_array(29)(142),
      output(30) => mem_array(30)(142),
      output(31) => mem_array(31)(142),
      output(32) => mem_array(32)(142),
      output(33) => mem_array(33)(142),
      output(34) => mem_array(34)(142),
      output(35) => mem_array(35)(142)
      );
  rom143 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001000000100000111100110000000000")
    port map (
      enable_o   => mem_enable_lines(143),
      output(0)  => mem_array(0)(143),
      output(1)  => mem_array(1)(143),
      output(2)  => mem_array(2)(143),
      output(3)  => mem_array(3)(143),
      output(4)  => mem_array(4)(143),
      output(5)  => mem_array(5)(143),
      output(6)  => mem_array(6)(143),
      output(7)  => mem_array(7)(143),
      output(8)  => mem_array(8)(143),
      output(9)  => mem_array(9)(143),
      output(10) => mem_array(10)(143),
      output(11) => mem_array(11)(143),
      output(12) => mem_array(12)(143),
      output(13) => mem_array(13)(143),
      output(14) => mem_array(14)(143),
      output(15) => mem_array(15)(143),
      output(16) => mem_array(16)(143),
      output(17) => mem_array(17)(143),
      output(18) => mem_array(18)(143),
      output(19) => mem_array(19)(143),
      output(20) => mem_array(20)(143),
      output(21) => mem_array(21)(143),
      output(22) => mem_array(22)(143),
      output(23) => mem_array(23)(143),
      output(24) => mem_array(24)(143),
      output(25) => mem_array(25)(143),
      output(26) => mem_array(26)(143),
      output(27) => mem_array(27)(143),
      output(28) => mem_array(28)(143),
      output(29) => mem_array(29)(143),
      output(30) => mem_array(30)(143),
      output(31) => mem_array(31)(143),
      output(32) => mem_array(32)(143),
      output(33) => mem_array(33)(143),
      output(34) => mem_array(34)(143),
      output(35) => mem_array(35)(143)
      );
  rom144 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000000100000100000011110011000000")
    port map (
      enable_o   => mem_enable_lines(144),
      output(0)  => mem_array(0)(144),
      output(1)  => mem_array(1)(144),
      output(2)  => mem_array(2)(144),
      output(3)  => mem_array(3)(144),
      output(4)  => mem_array(4)(144),
      output(5)  => mem_array(5)(144),
      output(6)  => mem_array(6)(144),
      output(7)  => mem_array(7)(144),
      output(8)  => mem_array(8)(144),
      output(9)  => mem_array(9)(144),
      output(10) => mem_array(10)(144),
      output(11) => mem_array(11)(144),
      output(12) => mem_array(12)(144),
      output(13) => mem_array(13)(144),
      output(14) => mem_array(14)(144),
      output(15) => mem_array(15)(144),
      output(16) => mem_array(16)(144),
      output(17) => mem_array(17)(144),
      output(18) => mem_array(18)(144),
      output(19) => mem_array(19)(144),
      output(20) => mem_array(20)(144),
      output(21) => mem_array(21)(144),
      output(22) => mem_array(22)(144),
      output(23) => mem_array(23)(144),
      output(24) => mem_array(24)(144),
      output(25) => mem_array(25)(144),
      output(26) => mem_array(26)(144),
      output(27) => mem_array(27)(144),
      output(28) => mem_array(28)(144),
      output(29) => mem_array(29)(144),
      output(30) => mem_array(30)(144),
      output(31) => mem_array(31)(144),
      output(32) => mem_array(32)(144),
      output(33) => mem_array(33)(144),
      output(34) => mem_array(34)(144),
      output(35) => mem_array(35)(144)
      );
  rom145 : entity work.rom
    generic map (
      bits  => 36,
      value => "000010000000010000011000001111011100")
    port map (
      enable_o   => mem_enable_lines(145),
      output(0)  => mem_array(0)(145),
      output(1)  => mem_array(1)(145),
      output(2)  => mem_array(2)(145),
      output(3)  => mem_array(3)(145),
      output(4)  => mem_array(4)(145),
      output(5)  => mem_array(5)(145),
      output(6)  => mem_array(6)(145),
      output(7)  => mem_array(7)(145),
      output(8)  => mem_array(8)(145),
      output(9)  => mem_array(9)(145),
      output(10) => mem_array(10)(145),
      output(11) => mem_array(11)(145),
      output(12) => mem_array(12)(145),
      output(13) => mem_array(13)(145),
      output(14) => mem_array(14)(145),
      output(15) => mem_array(15)(145),
      output(16) => mem_array(16)(145),
      output(17) => mem_array(17)(145),
      output(18) => mem_array(18)(145),
      output(19) => mem_array(19)(145),
      output(20) => mem_array(20)(145),
      output(21) => mem_array(21)(145),
      output(22) => mem_array(22)(145),
      output(23) => mem_array(23)(145),
      output(24) => mem_array(24)(145),
      output(25) => mem_array(25)(145),
      output(26) => mem_array(26)(145),
      output(27) => mem_array(27)(145),
      output(28) => mem_array(28)(145),
      output(29) => mem_array(29)(145),
      output(30) => mem_array(30)(145),
      output(31) => mem_array(31)(145),
      output(32) => mem_array(32)(145),
      output(33) => mem_array(33)(145),
      output(34) => mem_array(34)(145),
      output(35) => mem_array(35)(145)
      );
  rom146 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000001000000001000010100000111100")
    port map (
      enable_o   => mem_enable_lines(146),
      output(0)  => mem_array(0)(146),
      output(1)  => mem_array(1)(146),
      output(2)  => mem_array(2)(146),
      output(3)  => mem_array(3)(146),
      output(4)  => mem_array(4)(146),
      output(5)  => mem_array(5)(146),
      output(6)  => mem_array(6)(146),
      output(7)  => mem_array(7)(146),
      output(8)  => mem_array(8)(146),
      output(9)  => mem_array(9)(146),
      output(10) => mem_array(10)(146),
      output(11) => mem_array(11)(146),
      output(12) => mem_array(12)(146),
      output(13) => mem_array(13)(146),
      output(14) => mem_array(14)(146),
      output(15) => mem_array(15)(146),
      output(16) => mem_array(16)(146),
      output(17) => mem_array(17)(146),
      output(18) => mem_array(18)(146),
      output(19) => mem_array(19)(146),
      output(20) => mem_array(20)(146),
      output(21) => mem_array(21)(146),
      output(22) => mem_array(22)(146),
      output(23) => mem_array(23)(146),
      output(24) => mem_array(24)(146),
      output(25) => mem_array(25)(146),
      output(26) => mem_array(26)(146),
      output(27) => mem_array(27)(146),
      output(28) => mem_array(28)(146),
      output(29) => mem_array(29)(146),
      output(30) => mem_array(30)(146),
      output(31) => mem_array(31)(146),
      output(32) => mem_array(32)(146),
      output(33) => mem_array(33)(146),
      output(34) => mem_array(34)(146),
      output(35) => mem_array(35)(146)
      );
  rom147 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000010100100000000001010100000001")
    port map (
      enable_o   => mem_enable_lines(147),
      output(0)  => mem_array(0)(147),
      output(1)  => mem_array(1)(147),
      output(2)  => mem_array(2)(147),
      output(3)  => mem_array(3)(147),
      output(4)  => mem_array(4)(147),
      output(5)  => mem_array(5)(147),
      output(6)  => mem_array(6)(147),
      output(7)  => mem_array(7)(147),
      output(8)  => mem_array(8)(147),
      output(9)  => mem_array(9)(147),
      output(10) => mem_array(10)(147),
      output(11) => mem_array(11)(147),
      output(12) => mem_array(12)(147),
      output(13) => mem_array(13)(147),
      output(14) => mem_array(14)(147),
      output(15) => mem_array(15)(147),
      output(16) => mem_array(16)(147),
      output(17) => mem_array(17)(147),
      output(18) => mem_array(18)(147),
      output(19) => mem_array(19)(147),
      output(20) => mem_array(20)(147),
      output(21) => mem_array(21)(147),
      output(22) => mem_array(22)(147),
      output(23) => mem_array(23)(147),
      output(24) => mem_array(24)(147),
      output(25) => mem_array(25)(147),
      output(26) => mem_array(26)(147),
      output(27) => mem_array(27)(147),
      output(28) => mem_array(28)(147),
      output(29) => mem_array(29)(147),
      output(30) => mem_array(30)(147),
      output(31) => mem_array(31)(147),
      output(32) => mem_array(32)(147),
      output(33) => mem_array(33)(147),
      output(34) => mem_array(34)(147),
      output(35) => mem_array(35)(147)
      );
  rom148 : entity work.rom
    generic map (
      bits  => 36,
      value => "010010000000000001010000011111111000")
    port map (
      enable_o   => mem_enable_lines(148),
      output(0)  => mem_array(0)(148),
      output(1)  => mem_array(1)(148),
      output(2)  => mem_array(2)(148),
      output(3)  => mem_array(3)(148),
      output(4)  => mem_array(4)(148),
      output(5)  => mem_array(5)(148),
      output(6)  => mem_array(6)(148),
      output(7)  => mem_array(7)(148),
      output(8)  => mem_array(8)(148),
      output(9)  => mem_array(9)(148),
      output(10) => mem_array(10)(148),
      output(11) => mem_array(11)(148),
      output(12) => mem_array(12)(148),
      output(13) => mem_array(13)(148),
      output(14) => mem_array(14)(148),
      output(15) => mem_array(15)(148),
      output(16) => mem_array(16)(148),
      output(17) => mem_array(17)(148),
      output(18) => mem_array(18)(148),
      output(19) => mem_array(19)(148),
      output(20) => mem_array(20)(148),
      output(21) => mem_array(21)(148),
      output(22) => mem_array(22)(148),
      output(23) => mem_array(23)(148),
      output(24) => mem_array(24)(148),
      output(25) => mem_array(25)(148),
      output(26) => mem_array(26)(148),
      output(27) => mem_array(27)(148),
      output(28) => mem_array(28)(148),
      output(29) => mem_array(29)(148),
      output(30) => mem_array(30)(148),
      output(31) => mem_array(31)(148),
      output(32) => mem_array(32)(148),
      output(33) => mem_array(33)(148),
      output(34) => mem_array(34)(148),
      output(35) => mem_array(35)(148)
      );
  rom149 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001000011")
    port map (
      enable_o   => mem_enable_lines(149),
      output(0)  => mem_array(0)(149),
      output(1)  => mem_array(1)(149),
      output(2)  => mem_array(2)(149),
      output(3)  => mem_array(3)(149),
      output(4)  => mem_array(4)(149),
      output(5)  => mem_array(5)(149),
      output(6)  => mem_array(6)(149),
      output(7)  => mem_array(7)(149),
      output(8)  => mem_array(8)(149),
      output(9)  => mem_array(9)(149),
      output(10) => mem_array(10)(149),
      output(11) => mem_array(11)(149),
      output(12) => mem_array(12)(149),
      output(13) => mem_array(13)(149),
      output(14) => mem_array(14)(149),
      output(15) => mem_array(15)(149),
      output(16) => mem_array(16)(149),
      output(17) => mem_array(17)(149),
      output(18) => mem_array(18)(149),
      output(19) => mem_array(19)(149),
      output(20) => mem_array(20)(149),
      output(21) => mem_array(21)(149),
      output(22) => mem_array(22)(149),
      output(23) => mem_array(23)(149),
      output(24) => mem_array(24)(149),
      output(25) => mem_array(25)(149),
      output(26) => mem_array(26)(149),
      output(27) => mem_array(27)(149),
      output(28) => mem_array(28)(149),
      output(29) => mem_array(29)(149),
      output(30) => mem_array(30)(149),
      output(31) => mem_array(31)(149),
      output(32) => mem_array(32)(149),
      output(33) => mem_array(33)(149),
      output(34) => mem_array(34)(149),
      output(35) => mem_array(35)(149)
      );
  rom150 : entity work.rom
    generic map (
      bits  => 36,
      value => "100000111100010000000000100000000100")
    port map (
      enable_o   => mem_enable_lines(150),
      output(0)  => mem_array(0)(150),
      output(1)  => mem_array(1)(150),
      output(2)  => mem_array(2)(150),
      output(3)  => mem_array(3)(150),
      output(4)  => mem_array(4)(150),
      output(5)  => mem_array(5)(150),
      output(6)  => mem_array(6)(150),
      output(7)  => mem_array(7)(150),
      output(8)  => mem_array(8)(150),
      output(9)  => mem_array(9)(150),
      output(10) => mem_array(10)(150),
      output(11) => mem_array(11)(150),
      output(12) => mem_array(12)(150),
      output(13) => mem_array(13)(150),
      output(14) => mem_array(14)(150),
      output(15) => mem_array(15)(150),
      output(16) => mem_array(16)(150),
      output(17) => mem_array(17)(150),
      output(18) => mem_array(18)(150),
      output(19) => mem_array(19)(150),
      output(20) => mem_array(20)(150),
      output(21) => mem_array(21)(150),
      output(22) => mem_array(22)(150),
      output(23) => mem_array(23)(150),
      output(24) => mem_array(24)(150),
      output(25) => mem_array(25)(150),
      output(26) => mem_array(26)(150),
      output(27) => mem_array(27)(150),
      output(28) => mem_array(28)(150),
      output(29) => mem_array(29)(150),
      output(30) => mem_array(30)(150),
      output(31) => mem_array(31)(150),
      output(32) => mem_array(32)(150),
      output(33) => mem_array(33)(150),
      output(34) => mem_array(34)(150),
      output(35) => mem_array(35)(150)
      );
  rom151 : entity work.rom
    generic map (
      bits  => 36,
      value => "010000000011110000000000100010000000")
    port map (
      enable_o   => mem_enable_lines(151),
      output(0)  => mem_array(0)(151),
      output(1)  => mem_array(1)(151),
      output(2)  => mem_array(2)(151),
      output(3)  => mem_array(3)(151),
      output(4)  => mem_array(4)(151),
      output(5)  => mem_array(5)(151),
      output(6)  => mem_array(6)(151),
      output(7)  => mem_array(7)(151),
      output(8)  => mem_array(8)(151),
      output(9)  => mem_array(9)(151),
      output(10) => mem_array(10)(151),
      output(11) => mem_array(11)(151),
      output(12) => mem_array(12)(151),
      output(13) => mem_array(13)(151),
      output(14) => mem_array(14)(151),
      output(15) => mem_array(15)(151),
      output(16) => mem_array(16)(151),
      output(17) => mem_array(17)(151),
      output(18) => mem_array(18)(151),
      output(19) => mem_array(19)(151),
      output(20) => mem_array(20)(151),
      output(21) => mem_array(21)(151),
      output(22) => mem_array(22)(151),
      output(23) => mem_array(23)(151),
      output(24) => mem_array(24)(151),
      output(25) => mem_array(25)(151),
      output(26) => mem_array(26)(151),
      output(27) => mem_array(27)(151),
      output(28) => mem_array(28)(151),
      output(29) => mem_array(29)(151),
      output(30) => mem_array(30)(151),
      output(31) => mem_array(31)(151),
      output(32) => mem_array(32)(151),
      output(33) => mem_array(33)(151),
      output(34) => mem_array(34)(151),
      output(35) => mem_array(35)(151)
      );
  rom152 : entity work.rom
    generic map (
      bits  => 36,
      value => "010001001000000101000000000101000111")
    port map (
      enable_o   => mem_enable_lines(152),
      output(0)  => mem_array(0)(152),
      output(1)  => mem_array(1)(152),
      output(2)  => mem_array(2)(152),
      output(3)  => mem_array(3)(152),
      output(4)  => mem_array(4)(152),
      output(5)  => mem_array(5)(152),
      output(6)  => mem_array(6)(152),
      output(7)  => mem_array(7)(152),
      output(8)  => mem_array(8)(152),
      output(9)  => mem_array(9)(152),
      output(10) => mem_array(10)(152),
      output(11) => mem_array(11)(152),
      output(12) => mem_array(12)(152),
      output(13) => mem_array(13)(152),
      output(14) => mem_array(14)(152),
      output(15) => mem_array(15)(152),
      output(16) => mem_array(16)(152),
      output(17) => mem_array(17)(152),
      output(18) => mem_array(18)(152),
      output(19) => mem_array(19)(152),
      output(20) => mem_array(20)(152),
      output(21) => mem_array(21)(152),
      output(22) => mem_array(22)(152),
      output(23) => mem_array(23)(152),
      output(24) => mem_array(24)(152),
      output(25) => mem_array(25)(152),
      output(26) => mem_array(26)(152),
      output(27) => mem_array(27)(152),
      output(28) => mem_array(28)(152),
      output(29) => mem_array(29)(152),
      output(30) => mem_array(30)(152),
      output(31) => mem_array(31)(152),
      output(32) => mem_array(32)(152),
      output(33) => mem_array(33)(152),
      output(34) => mem_array(34)(152),
      output(35) => mem_array(35)(152)
      );
  rom153 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001000101000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(153),
      output(0)  => mem_array(0)(153),
      output(1)  => mem_array(1)(153),
      output(2)  => mem_array(2)(153),
      output(3)  => mem_array(3)(153),
      output(4)  => mem_array(4)(153),
      output(5)  => mem_array(5)(153),
      output(6)  => mem_array(6)(153),
      output(7)  => mem_array(7)(153),
      output(8)  => mem_array(8)(153),
      output(9)  => mem_array(9)(153),
      output(10) => mem_array(10)(153),
      output(11) => mem_array(11)(153),
      output(12) => mem_array(12)(153),
      output(13) => mem_array(13)(153),
      output(14) => mem_array(14)(153),
      output(15) => mem_array(15)(153),
      output(16) => mem_array(16)(153),
      output(17) => mem_array(17)(153),
      output(18) => mem_array(18)(153),
      output(19) => mem_array(19)(153),
      output(20) => mem_array(20)(153),
      output(21) => mem_array(21)(153),
      output(22) => mem_array(22)(153),
      output(23) => mem_array(23)(153),
      output(24) => mem_array(24)(153),
      output(25) => mem_array(25)(153),
      output(26) => mem_array(26)(153),
      output(27) => mem_array(27)(153),
      output(28) => mem_array(28)(153),
      output(29) => mem_array(29)(153),
      output(30) => mem_array(30)(153),
      output(31) => mem_array(31)(153),
      output(32) => mem_array(32)(153),
      output(33) => mem_array(33)(153),
      output(34) => mem_array(34)(153),
      output(35) => mem_array(35)(153)
      );
  rom154 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000100010110000011011000000100")
    port map (
      enable_o   => mem_enable_lines(154),
      output(0)  => mem_array(0)(154),
      output(1)  => mem_array(1)(154),
      output(2)  => mem_array(2)(154),
      output(3)  => mem_array(3)(154),
      output(4)  => mem_array(4)(154),
      output(5)  => mem_array(5)(154),
      output(6)  => mem_array(6)(154),
      output(7)  => mem_array(7)(154),
      output(8)  => mem_array(8)(154),
      output(9)  => mem_array(9)(154),
      output(10) => mem_array(10)(154),
      output(11) => mem_array(11)(154),
      output(12) => mem_array(12)(154),
      output(13) => mem_array(13)(154),
      output(14) => mem_array(14)(154),
      output(15) => mem_array(15)(154),
      output(16) => mem_array(16)(154),
      output(17) => mem_array(17)(154),
      output(18) => mem_array(18)(154),
      output(19) => mem_array(19)(154),
      output(20) => mem_array(20)(154),
      output(21) => mem_array(21)(154),
      output(22) => mem_array(22)(154),
      output(23) => mem_array(23)(154),
      output(24) => mem_array(24)(154),
      output(25) => mem_array(25)(154),
      output(26) => mem_array(26)(154),
      output(27) => mem_array(27)(154),
      output(28) => mem_array(28)(154),
      output(29) => mem_array(29)(154),
      output(30) => mem_array(30)(154),
      output(31) => mem_array(31)(154),
      output(32) => mem_array(32)(154),
      output(33) => mem_array(33)(154),
      output(34) => mem_array(34)(154),
      output(35) => mem_array(35)(154)
      );
  rom155 : entity work.rom
    generic map (
      bits  => 36,
      value => "101001000000010001100000000000000000")
    port map (
      enable_o   => mem_enable_lines(155),
      output(0)  => mem_array(0)(155),
      output(1)  => mem_array(1)(155),
      output(2)  => mem_array(2)(155),
      output(3)  => mem_array(3)(155),
      output(4)  => mem_array(4)(155),
      output(5)  => mem_array(5)(155),
      output(6)  => mem_array(6)(155),
      output(7)  => mem_array(7)(155),
      output(8)  => mem_array(8)(155),
      output(9)  => mem_array(9)(155),
      output(10) => mem_array(10)(155),
      output(11) => mem_array(11)(155),
      output(12) => mem_array(12)(155),
      output(13) => mem_array(13)(155),
      output(14) => mem_array(14)(155),
      output(15) => mem_array(15)(155),
      output(16) => mem_array(16)(155),
      output(17) => mem_array(17)(155),
      output(18) => mem_array(18)(155),
      output(19) => mem_array(19)(155),
      output(20) => mem_array(20)(155),
      output(21) => mem_array(21)(155),
      output(22) => mem_array(22)(155),
      output(23) => mem_array(23)(155),
      output(24) => mem_array(24)(155),
      output(25) => mem_array(25)(155),
      output(26) => mem_array(26)(155),
      output(27) => mem_array(27)(155),
      output(28) => mem_array(28)(155),
      output(29) => mem_array(29)(155),
      output(30) => mem_array(30)(155),
      output(31) => mem_array(31)(155),
      output(32) => mem_array(32)(155),
      output(33) => mem_array(33)(155),
      output(34) => mem_array(34)(155),
      output(35) => mem_array(35)(155)
      );
  rom156 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000001000000010100")
    port map (
      enable_o   => mem_enable_lines(156),
      output(0)  => mem_array(0)(156),
      output(1)  => mem_array(1)(156),
      output(2)  => mem_array(2)(156),
      output(3)  => mem_array(3)(156),
      output(4)  => mem_array(4)(156),
      output(5)  => mem_array(5)(156),
      output(6)  => mem_array(6)(156),
      output(7)  => mem_array(7)(156),
      output(8)  => mem_array(8)(156),
      output(9)  => mem_array(9)(156),
      output(10) => mem_array(10)(156),
      output(11) => mem_array(11)(156),
      output(12) => mem_array(12)(156),
      output(13) => mem_array(13)(156),
      output(14) => mem_array(14)(156),
      output(15) => mem_array(15)(156),
      output(16) => mem_array(16)(156),
      output(17) => mem_array(17)(156),
      output(18) => mem_array(18)(156),
      output(19) => mem_array(19)(156),
      output(20) => mem_array(20)(156),
      output(21) => mem_array(21)(156),
      output(22) => mem_array(22)(156),
      output(23) => mem_array(23)(156),
      output(24) => mem_array(24)(156),
      output(25) => mem_array(25)(156),
      output(26) => mem_array(26)(156),
      output(27) => mem_array(27)(156),
      output(28) => mem_array(28)(156),
      output(29) => mem_array(29)(156),
      output(30) => mem_array(30)(156),
      output(31) => mem_array(31)(156),
      output(32) => mem_array(32)(156),
      output(33) => mem_array(33)(156),
      output(34) => mem_array(34)(156),
      output(35) => mem_array(35)(156)
      );
  rom157 : entity work.rom
    generic map (
      bits  => 36,
      value => "001000000000000000000100011100000011")
    port map (
      enable_o   => mem_enable_lines(157),
      output(0)  => mem_array(0)(157),
      output(1)  => mem_array(1)(157),
      output(2)  => mem_array(2)(157),
      output(3)  => mem_array(3)(157),
      output(4)  => mem_array(4)(157),
      output(5)  => mem_array(5)(157),
      output(6)  => mem_array(6)(157),
      output(7)  => mem_array(7)(157),
      output(8)  => mem_array(8)(157),
      output(9)  => mem_array(9)(157),
      output(10) => mem_array(10)(157),
      output(11) => mem_array(11)(157),
      output(12) => mem_array(12)(157),
      output(13) => mem_array(13)(157),
      output(14) => mem_array(14)(157),
      output(15) => mem_array(15)(157),
      output(16) => mem_array(16)(157),
      output(17) => mem_array(17)(157),
      output(18) => mem_array(18)(157),
      output(19) => mem_array(19)(157),
      output(20) => mem_array(20)(157),
      output(21) => mem_array(21)(157),
      output(22) => mem_array(22)(157),
      output(23) => mem_array(23)(157),
      output(24) => mem_array(24)(157),
      output(25) => mem_array(25)(157),
      output(26) => mem_array(26)(157),
      output(27) => mem_array(27)(157),
      output(28) => mem_array(28)(157),
      output(29) => mem_array(29)(157),
      output(30) => mem_array(30)(157),
      output(31) => mem_array(31)(157),
      output(32) => mem_array(32)(157),
      output(33) => mem_array(33)(157),
      output(34) => mem_array(34)(157),
      output(35) => mem_array(35)(157)
      );
  rom158 : entity work.rom
    generic map (
      bits  => 36,
      value => "110001000000000010000000010001111000")
    port map (
      enable_o   => mem_enable_lines(158),
      output(0)  => mem_array(0)(158),
      output(1)  => mem_array(1)(158),
      output(2)  => mem_array(2)(158),
      output(3)  => mem_array(3)(158),
      output(4)  => mem_array(4)(158),
      output(5)  => mem_array(5)(158),
      output(6)  => mem_array(6)(158),
      output(7)  => mem_array(7)(158),
      output(8)  => mem_array(8)(158),
      output(9)  => mem_array(9)(158),
      output(10) => mem_array(10)(158),
      output(11) => mem_array(11)(158),
      output(12) => mem_array(12)(158),
      output(13) => mem_array(13)(158),
      output(14) => mem_array(14)(158),
      output(15) => mem_array(15)(158),
      output(16) => mem_array(16)(158),
      output(17) => mem_array(17)(158),
      output(18) => mem_array(18)(158),
      output(19) => mem_array(19)(158),
      output(20) => mem_array(20)(158),
      output(21) => mem_array(21)(158),
      output(22) => mem_array(22)(158),
      output(23) => mem_array(23)(158),
      output(24) => mem_array(24)(158),
      output(25) => mem_array(25)(158),
      output(26) => mem_array(26)(158),
      output(27) => mem_array(27)(158),
      output(28) => mem_array(28)(158),
      output(29) => mem_array(29)(158),
      output(30) => mem_array(30)(158),
      output(31) => mem_array(31)(158),
      output(32) => mem_array(32)(158),
      output(33) => mem_array(33)(158),
      output(34) => mem_array(34)(158),
      output(35) => mem_array(35)(158)
      );
  rom159 : entity work.rom
    generic map (
      bits  => 36,
      value => "001111000000000010101000000001001000")
    port map (
      enable_o   => mem_enable_lines(159),
      output(0)  => mem_array(0)(159),
      output(1)  => mem_array(1)(159),
      output(2)  => mem_array(2)(159),
      output(3)  => mem_array(3)(159),
      output(4)  => mem_array(4)(159),
      output(5)  => mem_array(5)(159),
      output(6)  => mem_array(6)(159),
      output(7)  => mem_array(7)(159),
      output(8)  => mem_array(8)(159),
      output(9)  => mem_array(9)(159),
      output(10) => mem_array(10)(159),
      output(11) => mem_array(11)(159),
      output(12) => mem_array(12)(159),
      output(13) => mem_array(13)(159),
      output(14) => mem_array(14)(159),
      output(15) => mem_array(15)(159),
      output(16) => mem_array(16)(159),
      output(17) => mem_array(17)(159),
      output(18) => mem_array(18)(159),
      output(19) => mem_array(19)(159),
      output(20) => mem_array(20)(159),
      output(21) => mem_array(21)(159),
      output(22) => mem_array(22)(159),
      output(23) => mem_array(23)(159),
      output(24) => mem_array(24)(159),
      output(25) => mem_array(25)(159),
      output(26) => mem_array(26)(159),
      output(27) => mem_array(27)(159),
      output(28) => mem_array(28)(159),
      output(29) => mem_array(29)(159),
      output(30) => mem_array(30)(159),
      output(31) => mem_array(31)(159),
      output(32) => mem_array(32)(159),
      output(33) => mem_array(33)(159),
      output(34) => mem_array(34)(159),
      output(35) => mem_array(35)(159)
      );
  rom160 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000110101000001001000010000000000")
    port map (
      enable_o   => mem_enable_lines(160),
      output(0)  => mem_array(0)(160),
      output(1)  => mem_array(1)(160),
      output(2)  => mem_array(2)(160),
      output(3)  => mem_array(3)(160),
      output(4)  => mem_array(4)(160),
      output(5)  => mem_array(5)(160),
      output(6)  => mem_array(6)(160),
      output(7)  => mem_array(7)(160),
      output(8)  => mem_array(8)(160),
      output(9)  => mem_array(9)(160),
      output(10) => mem_array(10)(160),
      output(11) => mem_array(11)(160),
      output(12) => mem_array(12)(160),
      output(13) => mem_array(13)(160),
      output(14) => mem_array(14)(160),
      output(15) => mem_array(15)(160),
      output(16) => mem_array(16)(160),
      output(17) => mem_array(17)(160),
      output(18) => mem_array(18)(160),
      output(19) => mem_array(19)(160),
      output(20) => mem_array(20)(160),
      output(21) => mem_array(21)(160),
      output(22) => mem_array(22)(160),
      output(23) => mem_array(23)(160),
      output(24) => mem_array(24)(160),
      output(25) => mem_array(25)(160),
      output(26) => mem_array(26)(160),
      output(27) => mem_array(27)(160),
      output(28) => mem_array(28)(160),
      output(29) => mem_array(29)(160),
      output(30) => mem_array(30)(160),
      output(31) => mem_array(31)(160),
      output(32) => mem_array(32)(160),
      output(33) => mem_array(33)(160),
      output(34) => mem_array(34)(160),
      output(35) => mem_array(35)(160)
      );
  rom161 : entity work.rom
    generic map (
      bits  => 36,
      value => "000100000001010000100000010000000000")
    port map (
      enable_o   => mem_enable_lines(161),
      output(0)  => mem_array(0)(161),
      output(1)  => mem_array(1)(161),
      output(2)  => mem_array(2)(161),
      output(3)  => mem_array(3)(161),
      output(4)  => mem_array(4)(161),
      output(5)  => mem_array(5)(161),
      output(6)  => mem_array(6)(161),
      output(7)  => mem_array(7)(161),
      output(8)  => mem_array(8)(161),
      output(9)  => mem_array(9)(161),
      output(10) => mem_array(10)(161),
      output(11) => mem_array(11)(161),
      output(12) => mem_array(12)(161),
      output(13) => mem_array(13)(161),
      output(14) => mem_array(14)(161),
      output(15) => mem_array(15)(161),
      output(16) => mem_array(16)(161),
      output(17) => mem_array(17)(161),
      output(18) => mem_array(18)(161),
      output(19) => mem_array(19)(161),
      output(20) => mem_array(20)(161),
      output(21) => mem_array(21)(161),
      output(22) => mem_array(22)(161),
      output(23) => mem_array(23)(161),
      output(24) => mem_array(24)(161),
      output(25) => mem_array(25)(161),
      output(26) => mem_array(26)(161),
      output(27) => mem_array(27)(161),
      output(28) => mem_array(28)(161),
      output(29) => mem_array(29)(161),
      output(30) => mem_array(30)(161),
      output(31) => mem_array(31)(161),
      output(32) => mem_array(32)(161),
      output(33) => mem_array(33)(161),
      output(34) => mem_array(34)(161),
      output(35) => mem_array(35)(161)
      );
  rom162 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(162),
      output(0)  => mem_array(0)(162),
      output(1)  => mem_array(1)(162),
      output(2)  => mem_array(2)(162),
      output(3)  => mem_array(3)(162),
      output(4)  => mem_array(4)(162),
      output(5)  => mem_array(5)(162),
      output(6)  => mem_array(6)(162),
      output(7)  => mem_array(7)(162),
      output(8)  => mem_array(8)(162),
      output(9)  => mem_array(9)(162),
      output(10) => mem_array(10)(162),
      output(11) => mem_array(11)(162),
      output(12) => mem_array(12)(162),
      output(13) => mem_array(13)(162),
      output(14) => mem_array(14)(162),
      output(15) => mem_array(15)(162),
      output(16) => mem_array(16)(162),
      output(17) => mem_array(17)(162),
      output(18) => mem_array(18)(162),
      output(19) => mem_array(19)(162),
      output(20) => mem_array(20)(162),
      output(21) => mem_array(21)(162),
      output(22) => mem_array(22)(162),
      output(23) => mem_array(23)(162),
      output(24) => mem_array(24)(162),
      output(25) => mem_array(25)(162),
      output(26) => mem_array(26)(162),
      output(27) => mem_array(27)(162),
      output(28) => mem_array(28)(162),
      output(29) => mem_array(29)(162),
      output(30) => mem_array(30)(162),
      output(31) => mem_array(31)(162),
      output(32) => mem_array(32)(162),
      output(33) => mem_array(33)(162),
      output(34) => mem_array(34)(162),
      output(35) => mem_array(35)(162)
      );
  rom163 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(163),
      output(0)  => mem_array(0)(163),
      output(1)  => mem_array(1)(163),
      output(2)  => mem_array(2)(163),
      output(3)  => mem_array(3)(163),
      output(4)  => mem_array(4)(163),
      output(5)  => mem_array(5)(163),
      output(6)  => mem_array(6)(163),
      output(7)  => mem_array(7)(163),
      output(8)  => mem_array(8)(163),
      output(9)  => mem_array(9)(163),
      output(10) => mem_array(10)(163),
      output(11) => mem_array(11)(163),
      output(12) => mem_array(12)(163),
      output(13) => mem_array(13)(163),
      output(14) => mem_array(14)(163),
      output(15) => mem_array(15)(163),
      output(16) => mem_array(16)(163),
      output(17) => mem_array(17)(163),
      output(18) => mem_array(18)(163),
      output(19) => mem_array(19)(163),
      output(20) => mem_array(20)(163),
      output(21) => mem_array(21)(163),
      output(22) => mem_array(22)(163),
      output(23) => mem_array(23)(163),
      output(24) => mem_array(24)(163),
      output(25) => mem_array(25)(163),
      output(26) => mem_array(26)(163),
      output(27) => mem_array(27)(163),
      output(28) => mem_array(28)(163),
      output(29) => mem_array(29)(163),
      output(30) => mem_array(30)(163),
      output(31) => mem_array(31)(163),
      output(32) => mem_array(32)(163),
      output(33) => mem_array(33)(163),
      output(34) => mem_array(34)(163),
      output(35) => mem_array(35)(163)
      );
  rom164 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(164),
      output(0)  => mem_array(0)(164),
      output(1)  => mem_array(1)(164),
      output(2)  => mem_array(2)(164),
      output(3)  => mem_array(3)(164),
      output(4)  => mem_array(4)(164),
      output(5)  => mem_array(5)(164),
      output(6)  => mem_array(6)(164),
      output(7)  => mem_array(7)(164),
      output(8)  => mem_array(8)(164),
      output(9)  => mem_array(9)(164),
      output(10) => mem_array(10)(164),
      output(11) => mem_array(11)(164),
      output(12) => mem_array(12)(164),
      output(13) => mem_array(13)(164),
      output(14) => mem_array(14)(164),
      output(15) => mem_array(15)(164),
      output(16) => mem_array(16)(164),
      output(17) => mem_array(17)(164),
      output(18) => mem_array(18)(164),
      output(19) => mem_array(19)(164),
      output(20) => mem_array(20)(164),
      output(21) => mem_array(21)(164),
      output(22) => mem_array(22)(164),
      output(23) => mem_array(23)(164),
      output(24) => mem_array(24)(164),
      output(25) => mem_array(25)(164),
      output(26) => mem_array(26)(164),
      output(27) => mem_array(27)(164),
      output(28) => mem_array(28)(164),
      output(29) => mem_array(29)(164),
      output(30) => mem_array(30)(164),
      output(31) => mem_array(31)(164),
      output(32) => mem_array(32)(164),
      output(33) => mem_array(33)(164),
      output(34) => mem_array(34)(164),
      output(35) => mem_array(35)(164)
      );
  rom165 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(165),
      output(0)  => mem_array(0)(165),
      output(1)  => mem_array(1)(165),
      output(2)  => mem_array(2)(165),
      output(3)  => mem_array(3)(165),
      output(4)  => mem_array(4)(165),
      output(5)  => mem_array(5)(165),
      output(6)  => mem_array(6)(165),
      output(7)  => mem_array(7)(165),
      output(8)  => mem_array(8)(165),
      output(9)  => mem_array(9)(165),
      output(10) => mem_array(10)(165),
      output(11) => mem_array(11)(165),
      output(12) => mem_array(12)(165),
      output(13) => mem_array(13)(165),
      output(14) => mem_array(14)(165),
      output(15) => mem_array(15)(165),
      output(16) => mem_array(16)(165),
      output(17) => mem_array(17)(165),
      output(18) => mem_array(18)(165),
      output(19) => mem_array(19)(165),
      output(20) => mem_array(20)(165),
      output(21) => mem_array(21)(165),
      output(22) => mem_array(22)(165),
      output(23) => mem_array(23)(165),
      output(24) => mem_array(24)(165),
      output(25) => mem_array(25)(165),
      output(26) => mem_array(26)(165),
      output(27) => mem_array(27)(165),
      output(28) => mem_array(28)(165),
      output(29) => mem_array(29)(165),
      output(30) => mem_array(30)(165),
      output(31) => mem_array(31)(165),
      output(32) => mem_array(32)(165),
      output(33) => mem_array(33)(165),
      output(34) => mem_array(34)(165),
      output(35) => mem_array(35)(165)
      );
  rom166 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(166),
      output(0)  => mem_array(0)(166),
      output(1)  => mem_array(1)(166),
      output(2)  => mem_array(2)(166),
      output(3)  => mem_array(3)(166),
      output(4)  => mem_array(4)(166),
      output(5)  => mem_array(5)(166),
      output(6)  => mem_array(6)(166),
      output(7)  => mem_array(7)(166),
      output(8)  => mem_array(8)(166),
      output(9)  => mem_array(9)(166),
      output(10) => mem_array(10)(166),
      output(11) => mem_array(11)(166),
      output(12) => mem_array(12)(166),
      output(13) => mem_array(13)(166),
      output(14) => mem_array(14)(166),
      output(15) => mem_array(15)(166),
      output(16) => mem_array(16)(166),
      output(17) => mem_array(17)(166),
      output(18) => mem_array(18)(166),
      output(19) => mem_array(19)(166),
      output(20) => mem_array(20)(166),
      output(21) => mem_array(21)(166),
      output(22) => mem_array(22)(166),
      output(23) => mem_array(23)(166),
      output(24) => mem_array(24)(166),
      output(25) => mem_array(25)(166),
      output(26) => mem_array(26)(166),
      output(27) => mem_array(27)(166),
      output(28) => mem_array(28)(166),
      output(29) => mem_array(29)(166),
      output(30) => mem_array(30)(166),
      output(31) => mem_array(31)(166),
      output(32) => mem_array(32)(166),
      output(33) => mem_array(33)(166),
      output(34) => mem_array(34)(166),
      output(35) => mem_array(35)(166)
      );
  rom167 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(167),
      output(0)  => mem_array(0)(167),
      output(1)  => mem_array(1)(167),
      output(2)  => mem_array(2)(167),
      output(3)  => mem_array(3)(167),
      output(4)  => mem_array(4)(167),
      output(5)  => mem_array(5)(167),
      output(6)  => mem_array(6)(167),
      output(7)  => mem_array(7)(167),
      output(8)  => mem_array(8)(167),
      output(9)  => mem_array(9)(167),
      output(10) => mem_array(10)(167),
      output(11) => mem_array(11)(167),
      output(12) => mem_array(12)(167),
      output(13) => mem_array(13)(167),
      output(14) => mem_array(14)(167),
      output(15) => mem_array(15)(167),
      output(16) => mem_array(16)(167),
      output(17) => mem_array(17)(167),
      output(18) => mem_array(18)(167),
      output(19) => mem_array(19)(167),
      output(20) => mem_array(20)(167),
      output(21) => mem_array(21)(167),
      output(22) => mem_array(22)(167),
      output(23) => mem_array(23)(167),
      output(24) => mem_array(24)(167),
      output(25) => mem_array(25)(167),
      output(26) => mem_array(26)(167),
      output(27) => mem_array(27)(167),
      output(28) => mem_array(28)(167),
      output(29) => mem_array(29)(167),
      output(30) => mem_array(30)(167),
      output(31) => mem_array(31)(167),
      output(32) => mem_array(32)(167),
      output(33) => mem_array(33)(167),
      output(34) => mem_array(34)(167),
      output(35) => mem_array(35)(167)
      );
  rom168 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(168),
      output(0)  => mem_array(0)(168),
      output(1)  => mem_array(1)(168),
      output(2)  => mem_array(2)(168),
      output(3)  => mem_array(3)(168),
      output(4)  => mem_array(4)(168),
      output(5)  => mem_array(5)(168),
      output(6)  => mem_array(6)(168),
      output(7)  => mem_array(7)(168),
      output(8)  => mem_array(8)(168),
      output(9)  => mem_array(9)(168),
      output(10) => mem_array(10)(168),
      output(11) => mem_array(11)(168),
      output(12) => mem_array(12)(168),
      output(13) => mem_array(13)(168),
      output(14) => mem_array(14)(168),
      output(15) => mem_array(15)(168),
      output(16) => mem_array(16)(168),
      output(17) => mem_array(17)(168),
      output(18) => mem_array(18)(168),
      output(19) => mem_array(19)(168),
      output(20) => mem_array(20)(168),
      output(21) => mem_array(21)(168),
      output(22) => mem_array(22)(168),
      output(23) => mem_array(23)(168),
      output(24) => mem_array(24)(168),
      output(25) => mem_array(25)(168),
      output(26) => mem_array(26)(168),
      output(27) => mem_array(27)(168),
      output(28) => mem_array(28)(168),
      output(29) => mem_array(29)(168),
      output(30) => mem_array(30)(168),
      output(31) => mem_array(31)(168),
      output(32) => mem_array(32)(168),
      output(33) => mem_array(33)(168),
      output(34) => mem_array(34)(168),
      output(35) => mem_array(35)(168)
      );
  rom169 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(169),
      output(0)  => mem_array(0)(169),
      output(1)  => mem_array(1)(169),
      output(2)  => mem_array(2)(169),
      output(3)  => mem_array(3)(169),
      output(4)  => mem_array(4)(169),
      output(5)  => mem_array(5)(169),
      output(6)  => mem_array(6)(169),
      output(7)  => mem_array(7)(169),
      output(8)  => mem_array(8)(169),
      output(9)  => mem_array(9)(169),
      output(10) => mem_array(10)(169),
      output(11) => mem_array(11)(169),
      output(12) => mem_array(12)(169),
      output(13) => mem_array(13)(169),
      output(14) => mem_array(14)(169),
      output(15) => mem_array(15)(169),
      output(16) => mem_array(16)(169),
      output(17) => mem_array(17)(169),
      output(18) => mem_array(18)(169),
      output(19) => mem_array(19)(169),
      output(20) => mem_array(20)(169),
      output(21) => mem_array(21)(169),
      output(22) => mem_array(22)(169),
      output(23) => mem_array(23)(169),
      output(24) => mem_array(24)(169),
      output(25) => mem_array(25)(169),
      output(26) => mem_array(26)(169),
      output(27) => mem_array(27)(169),
      output(28) => mem_array(28)(169),
      output(29) => mem_array(29)(169),
      output(30) => mem_array(30)(169),
      output(31) => mem_array(31)(169),
      output(32) => mem_array(32)(169),
      output(33) => mem_array(33)(169),
      output(34) => mem_array(34)(169),
      output(35) => mem_array(35)(169)
      );
  rom170 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000001")
    port map (
      enable_o   => mem_enable_lines(170),
      output(0)  => mem_array(0)(170),
      output(1)  => mem_array(1)(170),
      output(2)  => mem_array(2)(170),
      output(3)  => mem_array(3)(170),
      output(4)  => mem_array(4)(170),
      output(5)  => mem_array(5)(170),
      output(6)  => mem_array(6)(170),
      output(7)  => mem_array(7)(170),
      output(8)  => mem_array(8)(170),
      output(9)  => mem_array(9)(170),
      output(10) => mem_array(10)(170),
      output(11) => mem_array(11)(170),
      output(12) => mem_array(12)(170),
      output(13) => mem_array(13)(170),
      output(14) => mem_array(14)(170),
      output(15) => mem_array(15)(170),
      output(16) => mem_array(16)(170),
      output(17) => mem_array(17)(170),
      output(18) => mem_array(18)(170),
      output(19) => mem_array(19)(170),
      output(20) => mem_array(20)(170),
      output(21) => mem_array(21)(170),
      output(22) => mem_array(22)(170),
      output(23) => mem_array(23)(170),
      output(24) => mem_array(24)(170),
      output(25) => mem_array(25)(170),
      output(26) => mem_array(26)(170),
      output(27) => mem_array(27)(170),
      output(28) => mem_array(28)(170),
      output(29) => mem_array(29)(170),
      output(30) => mem_array(30)(170),
      output(31) => mem_array(31)(170),
      output(32) => mem_array(32)(170),
      output(33) => mem_array(33)(170),
      output(34) => mem_array(34)(170),
      output(35) => mem_array(35)(170)
      );
  rom171 : entity work.rom
    generic map (
      bits  => 36,
      value => "110000000011011000000100101001000000")
    port map (
      enable_o   => mem_enable_lines(171),
      output(0)  => mem_array(0)(171),
      output(1)  => mem_array(1)(171),
      output(2)  => mem_array(2)(171),
      output(3)  => mem_array(3)(171),
      output(4)  => mem_array(4)(171),
      output(5)  => mem_array(5)(171),
      output(6)  => mem_array(6)(171),
      output(7)  => mem_array(7)(171),
      output(8)  => mem_array(8)(171),
      output(9)  => mem_array(9)(171),
      output(10) => mem_array(10)(171),
      output(11) => mem_array(11)(171),
      output(12) => mem_array(12)(171),
      output(13) => mem_array(13)(171),
      output(14) => mem_array(14)(171),
      output(15) => mem_array(15)(171),
      output(16) => mem_array(16)(171),
      output(17) => mem_array(17)(171),
      output(18) => mem_array(18)(171),
      output(19) => mem_array(19)(171),
      output(20) => mem_array(20)(171),
      output(21) => mem_array(21)(171),
      output(22) => mem_array(22)(171),
      output(23) => mem_array(23)(171),
      output(24) => mem_array(24)(171),
      output(25) => mem_array(25)(171),
      output(26) => mem_array(26)(171),
      output(27) => mem_array(27)(171),
      output(28) => mem_array(28)(171),
      output(29) => mem_array(29)(171),
      output(30) => mem_array(30)(171),
      output(31) => mem_array(31)(171),
      output(32) => mem_array(32)(171),
      output(33) => mem_array(33)(171),
      output(34) => mem_array(34)(171),
      output(35) => mem_array(35)(171)
      );
  rom172 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(172),
      output(0)  => mem_array(0)(172),
      output(1)  => mem_array(1)(172),
      output(2)  => mem_array(2)(172),
      output(3)  => mem_array(3)(172),
      output(4)  => mem_array(4)(172),
      output(5)  => mem_array(5)(172),
      output(6)  => mem_array(6)(172),
      output(7)  => mem_array(7)(172),
      output(8)  => mem_array(8)(172),
      output(9)  => mem_array(9)(172),
      output(10) => mem_array(10)(172),
      output(11) => mem_array(11)(172),
      output(12) => mem_array(12)(172),
      output(13) => mem_array(13)(172),
      output(14) => mem_array(14)(172),
      output(15) => mem_array(15)(172),
      output(16) => mem_array(16)(172),
      output(17) => mem_array(17)(172),
      output(18) => mem_array(18)(172),
      output(19) => mem_array(19)(172),
      output(20) => mem_array(20)(172),
      output(21) => mem_array(21)(172),
      output(22) => mem_array(22)(172),
      output(23) => mem_array(23)(172),
      output(24) => mem_array(24)(172),
      output(25) => mem_array(25)(172),
      output(26) => mem_array(26)(172),
      output(27) => mem_array(27)(172),
      output(28) => mem_array(28)(172),
      output(29) => mem_array(29)(172),
      output(30) => mem_array(30)(172),
      output(31) => mem_array(31)(172),
      output(32) => mem_array(32)(172),
      output(33) => mem_array(33)(172),
      output(34) => mem_array(34)(172),
      output(35) => mem_array(35)(172)
      );
  rom173 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000011010000000110110000001001010")
    port map (
      enable_o   => mem_enable_lines(173),
      output(0)  => mem_array(0)(173),
      output(1)  => mem_array(1)(173),
      output(2)  => mem_array(2)(173),
      output(3)  => mem_array(3)(173),
      output(4)  => mem_array(4)(173),
      output(5)  => mem_array(5)(173),
      output(6)  => mem_array(6)(173),
      output(7)  => mem_array(7)(173),
      output(8)  => mem_array(8)(173),
      output(9)  => mem_array(9)(173),
      output(10) => mem_array(10)(173),
      output(11) => mem_array(11)(173),
      output(12) => mem_array(12)(173),
      output(13) => mem_array(13)(173),
      output(14) => mem_array(14)(173),
      output(15) => mem_array(15)(173),
      output(16) => mem_array(16)(173),
      output(17) => mem_array(17)(173),
      output(18) => mem_array(18)(173),
      output(19) => mem_array(19)(173),
      output(20) => mem_array(20)(173),
      output(21) => mem_array(21)(173),
      output(22) => mem_array(22)(173),
      output(23) => mem_array(23)(173),
      output(24) => mem_array(24)(173),
      output(25) => mem_array(25)(173),
      output(26) => mem_array(26)(173),
      output(27) => mem_array(27)(173),
      output(28) => mem_array(28)(173),
      output(29) => mem_array(29)(173),
      output(30) => mem_array(30)(173),
      output(31) => mem_array(31)(173),
      output(32) => mem_array(32)(173),
      output(33) => mem_array(33)(173),
      output(34) => mem_array(34)(173),
      output(35) => mem_array(35)(173)
      );
  rom174 : entity work.rom
    generic map (
      bits  => 36,
      value => "010000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(174),
      output(0)  => mem_array(0)(174),
      output(1)  => mem_array(1)(174),
      output(2)  => mem_array(2)(174),
      output(3)  => mem_array(3)(174),
      output(4)  => mem_array(4)(174),
      output(5)  => mem_array(5)(174),
      output(6)  => mem_array(6)(174),
      output(7)  => mem_array(7)(174),
      output(8)  => mem_array(8)(174),
      output(9)  => mem_array(9)(174),
      output(10) => mem_array(10)(174),
      output(11) => mem_array(11)(174),
      output(12) => mem_array(12)(174),
      output(13) => mem_array(13)(174),
      output(14) => mem_array(14)(174),
      output(15) => mem_array(15)(174),
      output(16) => mem_array(16)(174),
      output(17) => mem_array(17)(174),
      output(18) => mem_array(18)(174),
      output(19) => mem_array(19)(174),
      output(20) => mem_array(20)(174),
      output(21) => mem_array(21)(174),
      output(22) => mem_array(22)(174),
      output(23) => mem_array(23)(174),
      output(24) => mem_array(24)(174),
      output(25) => mem_array(25)(174),
      output(26) => mem_array(26)(174),
      output(27) => mem_array(27)(174),
      output(28) => mem_array(28)(174),
      output(29) => mem_array(29)(174),
      output(30) => mem_array(30)(174),
      output(31) => mem_array(31)(174),
      output(32) => mem_array(32)(174),
      output(33) => mem_array(33)(174),
      output(34) => mem_array(34)(174),
      output(35) => mem_array(35)(174)
      );
  rom175 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(175),
      output(0)  => mem_array(0)(175),
      output(1)  => mem_array(1)(175),
      output(2)  => mem_array(2)(175),
      output(3)  => mem_array(3)(175),
      output(4)  => mem_array(4)(175),
      output(5)  => mem_array(5)(175),
      output(6)  => mem_array(6)(175),
      output(7)  => mem_array(7)(175),
      output(8)  => mem_array(8)(175),
      output(9)  => mem_array(9)(175),
      output(10) => mem_array(10)(175),
      output(11) => mem_array(11)(175),
      output(12) => mem_array(12)(175),
      output(13) => mem_array(13)(175),
      output(14) => mem_array(14)(175),
      output(15) => mem_array(15)(175),
      output(16) => mem_array(16)(175),
      output(17) => mem_array(17)(175),
      output(18) => mem_array(18)(175),
      output(19) => mem_array(19)(175),
      output(20) => mem_array(20)(175),
      output(21) => mem_array(21)(175),
      output(22) => mem_array(22)(175),
      output(23) => mem_array(23)(175),
      output(24) => mem_array(24)(175),
      output(25) => mem_array(25)(175),
      output(26) => mem_array(26)(175),
      output(27) => mem_array(27)(175),
      output(28) => mem_array(28)(175),
      output(29) => mem_array(29)(175),
      output(30) => mem_array(30)(175),
      output(31) => mem_array(31)(175),
      output(32) => mem_array(32)(175),
      output(33) => mem_array(33)(175),
      output(34) => mem_array(34)(175),
      output(35) => mem_array(35)(175)
      );
  rom176 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(176),
      output(0)  => mem_array(0)(176),
      output(1)  => mem_array(1)(176),
      output(2)  => mem_array(2)(176),
      output(3)  => mem_array(3)(176),
      output(4)  => mem_array(4)(176),
      output(5)  => mem_array(5)(176),
      output(6)  => mem_array(6)(176),
      output(7)  => mem_array(7)(176),
      output(8)  => mem_array(8)(176),
      output(9)  => mem_array(9)(176),
      output(10) => mem_array(10)(176),
      output(11) => mem_array(11)(176),
      output(12) => mem_array(12)(176),
      output(13) => mem_array(13)(176),
      output(14) => mem_array(14)(176),
      output(15) => mem_array(15)(176),
      output(16) => mem_array(16)(176),
      output(17) => mem_array(17)(176),
      output(18) => mem_array(18)(176),
      output(19) => mem_array(19)(176),
      output(20) => mem_array(20)(176),
      output(21) => mem_array(21)(176),
      output(22) => mem_array(22)(176),
      output(23) => mem_array(23)(176),
      output(24) => mem_array(24)(176),
      output(25) => mem_array(25)(176),
      output(26) => mem_array(26)(176),
      output(27) => mem_array(27)(176),
      output(28) => mem_array(28)(176),
      output(29) => mem_array(29)(176),
      output(30) => mem_array(30)(176),
      output(31) => mem_array(31)(176),
      output(32) => mem_array(32)(176),
      output(33) => mem_array(33)(176),
      output(34) => mem_array(34)(176),
      output(35) => mem_array(35)(176)
      );
  rom177 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000001110110000011")
    port map (
      enable_o   => mem_enable_lines(177),
      output(0)  => mem_array(0)(177),
      output(1)  => mem_array(1)(177),
      output(2)  => mem_array(2)(177),
      output(3)  => mem_array(3)(177),
      output(4)  => mem_array(4)(177),
      output(5)  => mem_array(5)(177),
      output(6)  => mem_array(6)(177),
      output(7)  => mem_array(7)(177),
      output(8)  => mem_array(8)(177),
      output(9)  => mem_array(9)(177),
      output(10) => mem_array(10)(177),
      output(11) => mem_array(11)(177),
      output(12) => mem_array(12)(177),
      output(13) => mem_array(13)(177),
      output(14) => mem_array(14)(177),
      output(15) => mem_array(15)(177),
      output(16) => mem_array(16)(177),
      output(17) => mem_array(17)(177),
      output(18) => mem_array(18)(177),
      output(19) => mem_array(19)(177),
      output(20) => mem_array(20)(177),
      output(21) => mem_array(21)(177),
      output(22) => mem_array(22)(177),
      output(23) => mem_array(23)(177),
      output(24) => mem_array(24)(177),
      output(25) => mem_array(25)(177),
      output(26) => mem_array(26)(177),
      output(27) => mem_array(27)(177),
      output(28) => mem_array(28)(177),
      output(29) => mem_array(29)(177),
      output(30) => mem_array(30)(177),
      output(31) => mem_array(31)(177),
      output(32) => mem_array(32)(177),
      output(33) => mem_array(33)(177),
      output(34) => mem_array(34)(177),
      output(35) => mem_array(35)(177)
      );
  rom178 : entity work.rom
    generic map (
      bits  => 36,
      value => "011000000100101001000000011111110000")
    port map (
      enable_o   => mem_enable_lines(178),
      output(0)  => mem_array(0)(178),
      output(1)  => mem_array(1)(178),
      output(2)  => mem_array(2)(178),
      output(3)  => mem_array(3)(178),
      output(4)  => mem_array(4)(178),
      output(5)  => mem_array(5)(178),
      output(6)  => mem_array(6)(178),
      output(7)  => mem_array(7)(178),
      output(8)  => mem_array(8)(178),
      output(9)  => mem_array(9)(178),
      output(10) => mem_array(10)(178),
      output(11) => mem_array(11)(178),
      output(12) => mem_array(12)(178),
      output(13) => mem_array(13)(178),
      output(14) => mem_array(14)(178),
      output(15) => mem_array(15)(178),
      output(16) => mem_array(16)(178),
      output(17) => mem_array(17)(178),
      output(18) => mem_array(18)(178),
      output(19) => mem_array(19)(178),
      output(20) => mem_array(20)(178),
      output(21) => mem_array(21)(178),
      output(22) => mem_array(22)(178),
      output(23) => mem_array(23)(178),
      output(24) => mem_array(24)(178),
      output(25) => mem_array(25)(178),
      output(26) => mem_array(26)(178),
      output(27) => mem_array(27)(178),
      output(28) => mem_array(28)(178),
      output(29) => mem_array(29)(178),
      output(30) => mem_array(30)(178),
      output(31) => mem_array(31)(178),
      output(32) => mem_array(32)(178),
      output(33) => mem_array(33)(178),
      output(34) => mem_array(34)(178),
      output(35) => mem_array(35)(178)
      );
  rom179 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(179),
      output(0)  => mem_array(0)(179),
      output(1)  => mem_array(1)(179),
      output(2)  => mem_array(2)(179),
      output(3)  => mem_array(3)(179),
      output(4)  => mem_array(4)(179),
      output(5)  => mem_array(5)(179),
      output(6)  => mem_array(6)(179),
      output(7)  => mem_array(7)(179),
      output(8)  => mem_array(8)(179),
      output(9)  => mem_array(9)(179),
      output(10) => mem_array(10)(179),
      output(11) => mem_array(11)(179),
      output(12) => mem_array(12)(179),
      output(13) => mem_array(13)(179),
      output(14) => mem_array(14)(179),
      output(15) => mem_array(15)(179),
      output(16) => mem_array(16)(179),
      output(17) => mem_array(17)(179),
      output(18) => mem_array(18)(179),
      output(19) => mem_array(19)(179),
      output(20) => mem_array(20)(179),
      output(21) => mem_array(21)(179),
      output(22) => mem_array(22)(179),
      output(23) => mem_array(23)(179),
      output(24) => mem_array(24)(179),
      output(25) => mem_array(25)(179),
      output(26) => mem_array(26)(179),
      output(27) => mem_array(27)(179),
      output(28) => mem_array(28)(179),
      output(29) => mem_array(29)(179),
      output(30) => mem_array(30)(179),
      output(31) => mem_array(31)(179),
      output(32) => mem_array(32)(179),
      output(33) => mem_array(33)(179),
      output(34) => mem_array(34)(179),
      output(35) => mem_array(35)(179)
      );
  rom180 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(180),
      output(0)  => mem_array(0)(180),
      output(1)  => mem_array(1)(180),
      output(2)  => mem_array(2)(180),
      output(3)  => mem_array(3)(180),
      output(4)  => mem_array(4)(180),
      output(5)  => mem_array(5)(180),
      output(6)  => mem_array(6)(180),
      output(7)  => mem_array(7)(180),
      output(8)  => mem_array(8)(180),
      output(9)  => mem_array(9)(180),
      output(10) => mem_array(10)(180),
      output(11) => mem_array(11)(180),
      output(12) => mem_array(12)(180),
      output(13) => mem_array(13)(180),
      output(14) => mem_array(14)(180),
      output(15) => mem_array(15)(180),
      output(16) => mem_array(16)(180),
      output(17) => mem_array(17)(180),
      output(18) => mem_array(18)(180),
      output(19) => mem_array(19)(180),
      output(20) => mem_array(20)(180),
      output(21) => mem_array(21)(180),
      output(22) => mem_array(22)(180),
      output(23) => mem_array(23)(180),
      output(24) => mem_array(24)(180),
      output(25) => mem_array(25)(180),
      output(26) => mem_array(26)(180),
      output(27) => mem_array(27)(180),
      output(28) => mem_array(28)(180),
      output(29) => mem_array(29)(180),
      output(30) => mem_array(30)(180),
      output(31) => mem_array(31)(180),
      output(32) => mem_array(32)(180),
      output(33) => mem_array(33)(180),
      output(34) => mem_array(34)(180),
      output(35) => mem_array(35)(180)
      );
  rom181 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(181),
      output(0)  => mem_array(0)(181),
      output(1)  => mem_array(1)(181),
      output(2)  => mem_array(2)(181),
      output(3)  => mem_array(3)(181),
      output(4)  => mem_array(4)(181),
      output(5)  => mem_array(5)(181),
      output(6)  => mem_array(6)(181),
      output(7)  => mem_array(7)(181),
      output(8)  => mem_array(8)(181),
      output(9)  => mem_array(9)(181),
      output(10) => mem_array(10)(181),
      output(11) => mem_array(11)(181),
      output(12) => mem_array(12)(181),
      output(13) => mem_array(13)(181),
      output(14) => mem_array(14)(181),
      output(15) => mem_array(15)(181),
      output(16) => mem_array(16)(181),
      output(17) => mem_array(17)(181),
      output(18) => mem_array(18)(181),
      output(19) => mem_array(19)(181),
      output(20) => mem_array(20)(181),
      output(21) => mem_array(21)(181),
      output(22) => mem_array(22)(181),
      output(23) => mem_array(23)(181),
      output(24) => mem_array(24)(181),
      output(25) => mem_array(25)(181),
      output(26) => mem_array(26)(181),
      output(27) => mem_array(27)(181),
      output(28) => mem_array(28)(181),
      output(29) => mem_array(29)(181),
      output(30) => mem_array(30)(181),
      output(31) => mem_array(31)(181),
      output(32) => mem_array(32)(181),
      output(33) => mem_array(33)(181),
      output(34) => mem_array(34)(181),
      output(35) => mem_array(35)(181)
      );
  rom182 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(182),
      output(0)  => mem_array(0)(182),
      output(1)  => mem_array(1)(182),
      output(2)  => mem_array(2)(182),
      output(3)  => mem_array(3)(182),
      output(4)  => mem_array(4)(182),
      output(5)  => mem_array(5)(182),
      output(6)  => mem_array(6)(182),
      output(7)  => mem_array(7)(182),
      output(8)  => mem_array(8)(182),
      output(9)  => mem_array(9)(182),
      output(10) => mem_array(10)(182),
      output(11) => mem_array(11)(182),
      output(12) => mem_array(12)(182),
      output(13) => mem_array(13)(182),
      output(14) => mem_array(14)(182),
      output(15) => mem_array(15)(182),
      output(16) => mem_array(16)(182),
      output(17) => mem_array(17)(182),
      output(18) => mem_array(18)(182),
      output(19) => mem_array(19)(182),
      output(20) => mem_array(20)(182),
      output(21) => mem_array(21)(182),
      output(22) => mem_array(22)(182),
      output(23) => mem_array(23)(182),
      output(24) => mem_array(24)(182),
      output(25) => mem_array(25)(182),
      output(26) => mem_array(26)(182),
      output(27) => mem_array(27)(182),
      output(28) => mem_array(28)(182),
      output(29) => mem_array(29)(182),
      output(30) => mem_array(30)(182),
      output(31) => mem_array(31)(182),
      output(32) => mem_array(32)(182),
      output(33) => mem_array(33)(182),
      output(34) => mem_array(34)(182),
      output(35) => mem_array(35)(182)
      );
  rom183 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(183),
      output(0)  => mem_array(0)(183),
      output(1)  => mem_array(1)(183),
      output(2)  => mem_array(2)(183),
      output(3)  => mem_array(3)(183),
      output(4)  => mem_array(4)(183),
      output(5)  => mem_array(5)(183),
      output(6)  => mem_array(6)(183),
      output(7)  => mem_array(7)(183),
      output(8)  => mem_array(8)(183),
      output(9)  => mem_array(9)(183),
      output(10) => mem_array(10)(183),
      output(11) => mem_array(11)(183),
      output(12) => mem_array(12)(183),
      output(13) => mem_array(13)(183),
      output(14) => mem_array(14)(183),
      output(15) => mem_array(15)(183),
      output(16) => mem_array(16)(183),
      output(17) => mem_array(17)(183),
      output(18) => mem_array(18)(183),
      output(19) => mem_array(19)(183),
      output(20) => mem_array(20)(183),
      output(21) => mem_array(21)(183),
      output(22) => mem_array(22)(183),
      output(23) => mem_array(23)(183),
      output(24) => mem_array(24)(183),
      output(25) => mem_array(25)(183),
      output(26) => mem_array(26)(183),
      output(27) => mem_array(27)(183),
      output(28) => mem_array(28)(183),
      output(29) => mem_array(29)(183),
      output(30) => mem_array(30)(183),
      output(31) => mem_array(31)(183),
      output(32) => mem_array(32)(183),
      output(33) => mem_array(33)(183),
      output(34) => mem_array(34)(183),
      output(35) => mem_array(35)(183)
      );
  rom184 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(184),
      output(0)  => mem_array(0)(184),
      output(1)  => mem_array(1)(184),
      output(2)  => mem_array(2)(184),
      output(3)  => mem_array(3)(184),
      output(4)  => mem_array(4)(184),
      output(5)  => mem_array(5)(184),
      output(6)  => mem_array(6)(184),
      output(7)  => mem_array(7)(184),
      output(8)  => mem_array(8)(184),
      output(9)  => mem_array(9)(184),
      output(10) => mem_array(10)(184),
      output(11) => mem_array(11)(184),
      output(12) => mem_array(12)(184),
      output(13) => mem_array(13)(184),
      output(14) => mem_array(14)(184),
      output(15) => mem_array(15)(184),
      output(16) => mem_array(16)(184),
      output(17) => mem_array(17)(184),
      output(18) => mem_array(18)(184),
      output(19) => mem_array(19)(184),
      output(20) => mem_array(20)(184),
      output(21) => mem_array(21)(184),
      output(22) => mem_array(22)(184),
      output(23) => mem_array(23)(184),
      output(24) => mem_array(24)(184),
      output(25) => mem_array(25)(184),
      output(26) => mem_array(26)(184),
      output(27) => mem_array(27)(184),
      output(28) => mem_array(28)(184),
      output(29) => mem_array(29)(184),
      output(30) => mem_array(30)(184),
      output(31) => mem_array(31)(184),
      output(32) => mem_array(32)(184),
      output(33) => mem_array(33)(184),
      output(34) => mem_array(34)(184),
      output(35) => mem_array(35)(184)
      );
  rom185 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(185),
      output(0)  => mem_array(0)(185),
      output(1)  => mem_array(1)(185),
      output(2)  => mem_array(2)(185),
      output(3)  => mem_array(3)(185),
      output(4)  => mem_array(4)(185),
      output(5)  => mem_array(5)(185),
      output(6)  => mem_array(6)(185),
      output(7)  => mem_array(7)(185),
      output(8)  => mem_array(8)(185),
      output(9)  => mem_array(9)(185),
      output(10) => mem_array(10)(185),
      output(11) => mem_array(11)(185),
      output(12) => mem_array(12)(185),
      output(13) => mem_array(13)(185),
      output(14) => mem_array(14)(185),
      output(15) => mem_array(15)(185),
      output(16) => mem_array(16)(185),
      output(17) => mem_array(17)(185),
      output(18) => mem_array(18)(185),
      output(19) => mem_array(19)(185),
      output(20) => mem_array(20)(185),
      output(21) => mem_array(21)(185),
      output(22) => mem_array(22)(185),
      output(23) => mem_array(23)(185),
      output(24) => mem_array(24)(185),
      output(25) => mem_array(25)(185),
      output(26) => mem_array(26)(185),
      output(27) => mem_array(27)(185),
      output(28) => mem_array(28)(185),
      output(29) => mem_array(29)(185),
      output(30) => mem_array(30)(185),
      output(31) => mem_array(31)(185),
      output(32) => mem_array(32)(185),
      output(33) => mem_array(33)(185),
      output(34) => mem_array(34)(185),
      output(35) => mem_array(35)(185)
      );
  rom186 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000010111100000110110")
    port map (
      enable_o   => mem_enable_lines(186),
      output(0)  => mem_array(0)(186),
      output(1)  => mem_array(1)(186),
      output(2)  => mem_array(2)(186),
      output(3)  => mem_array(3)(186),
      output(4)  => mem_array(4)(186),
      output(5)  => mem_array(5)(186),
      output(6)  => mem_array(6)(186),
      output(7)  => mem_array(7)(186),
      output(8)  => mem_array(8)(186),
      output(9)  => mem_array(9)(186),
      output(10) => mem_array(10)(186),
      output(11) => mem_array(11)(186),
      output(12) => mem_array(12)(186),
      output(13) => mem_array(13)(186),
      output(14) => mem_array(14)(186),
      output(15) => mem_array(15)(186),
      output(16) => mem_array(16)(186),
      output(17) => mem_array(17)(186),
      output(18) => mem_array(18)(186),
      output(19) => mem_array(19)(186),
      output(20) => mem_array(20)(186),
      output(21) => mem_array(21)(186),
      output(22) => mem_array(22)(186),
      output(23) => mem_array(23)(186),
      output(24) => mem_array(24)(186),
      output(25) => mem_array(25)(186),
      output(26) => mem_array(26)(186),
      output(27) => mem_array(27)(186),
      output(28) => mem_array(28)(186),
      output(29) => mem_array(29)(186),
      output(30) => mem_array(30)(186),
      output(31) => mem_array(31)(186),
      output(32) => mem_array(32)(186),
      output(33) => mem_array(33)(186),
      output(34) => mem_array(34)(186),
      output(35) => mem_array(35)(186)
      );
  rom187 : entity work.rom
    generic map (
      bits  => 36,
      value => "010000000000000100000111111100000000")
    port map (
      enable_o   => mem_enable_lines(187),
      output(0)  => mem_array(0)(187),
      output(1)  => mem_array(1)(187),
      output(2)  => mem_array(2)(187),
      output(3)  => mem_array(3)(187),
      output(4)  => mem_array(4)(187),
      output(5)  => mem_array(5)(187),
      output(6)  => mem_array(6)(187),
      output(7)  => mem_array(7)(187),
      output(8)  => mem_array(8)(187),
      output(9)  => mem_array(9)(187),
      output(10) => mem_array(10)(187),
      output(11) => mem_array(11)(187),
      output(12) => mem_array(12)(187),
      output(13) => mem_array(13)(187),
      output(14) => mem_array(14)(187),
      output(15) => mem_array(15)(187),
      output(16) => mem_array(16)(187),
      output(17) => mem_array(17)(187),
      output(18) => mem_array(18)(187),
      output(19) => mem_array(19)(187),
      output(20) => mem_array(20)(187),
      output(21) => mem_array(21)(187),
      output(22) => mem_array(22)(187),
      output(23) => mem_array(23)(187),
      output(24) => mem_array(24)(187),
      output(25) => mem_array(25)(187),
      output(26) => mem_array(26)(187),
      output(27) => mem_array(27)(187),
      output(28) => mem_array(28)(187),
      output(29) => mem_array(29)(187),
      output(30) => mem_array(30)(187),
      output(31) => mem_array(31)(187),
      output(32) => mem_array(32)(187),
      output(33) => mem_array(33)(187),
      output(34) => mem_array(34)(187),
      output(35) => mem_array(35)(187)
      );
  rom188 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(188),
      output(0)  => mem_array(0)(188),
      output(1)  => mem_array(1)(188),
      output(2)  => mem_array(2)(188),
      output(3)  => mem_array(3)(188),
      output(4)  => mem_array(4)(188),
      output(5)  => mem_array(5)(188),
      output(6)  => mem_array(6)(188),
      output(7)  => mem_array(7)(188),
      output(8)  => mem_array(8)(188),
      output(9)  => mem_array(9)(188),
      output(10) => mem_array(10)(188),
      output(11) => mem_array(11)(188),
      output(12) => mem_array(12)(188),
      output(13) => mem_array(13)(188),
      output(14) => mem_array(14)(188),
      output(15) => mem_array(15)(188),
      output(16) => mem_array(16)(188),
      output(17) => mem_array(17)(188),
      output(18) => mem_array(18)(188),
      output(19) => mem_array(19)(188),
      output(20) => mem_array(20)(188),
      output(21) => mem_array(21)(188),
      output(22) => mem_array(22)(188),
      output(23) => mem_array(23)(188),
      output(24) => mem_array(24)(188),
      output(25) => mem_array(25)(188),
      output(26) => mem_array(26)(188),
      output(27) => mem_array(27)(188),
      output(28) => mem_array(28)(188),
      output(29) => mem_array(29)(188),
      output(30) => mem_array(30)(188),
      output(31) => mem_array(31)(188),
      output(32) => mem_array(32)(188),
      output(33) => mem_array(33)(188),
      output(34) => mem_array(34)(188),
      output(35) => mem_array(35)(188)
      );
  rom189 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(189),
      output(0)  => mem_array(0)(189),
      output(1)  => mem_array(1)(189),
      output(2)  => mem_array(2)(189),
      output(3)  => mem_array(3)(189),
      output(4)  => mem_array(4)(189),
      output(5)  => mem_array(5)(189),
      output(6)  => mem_array(6)(189),
      output(7)  => mem_array(7)(189),
      output(8)  => mem_array(8)(189),
      output(9)  => mem_array(9)(189),
      output(10) => mem_array(10)(189),
      output(11) => mem_array(11)(189),
      output(12) => mem_array(12)(189),
      output(13) => mem_array(13)(189),
      output(14) => mem_array(14)(189),
      output(15) => mem_array(15)(189),
      output(16) => mem_array(16)(189),
      output(17) => mem_array(17)(189),
      output(18) => mem_array(18)(189),
      output(19) => mem_array(19)(189),
      output(20) => mem_array(20)(189),
      output(21) => mem_array(21)(189),
      output(22) => mem_array(22)(189),
      output(23) => mem_array(23)(189),
      output(24) => mem_array(24)(189),
      output(25) => mem_array(25)(189),
      output(26) => mem_array(26)(189),
      output(27) => mem_array(27)(189),
      output(28) => mem_array(28)(189),
      output(29) => mem_array(29)(189),
      output(30) => mem_array(30)(189),
      output(31) => mem_array(31)(189),
      output(32) => mem_array(32)(189),
      output(33) => mem_array(33)(189),
      output(34) => mem_array(34)(189),
      output(35) => mem_array(35)(189)
      );
  rom190 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(190),
      output(0)  => mem_array(0)(190),
      output(1)  => mem_array(1)(190),
      output(2)  => mem_array(2)(190),
      output(3)  => mem_array(3)(190),
      output(4)  => mem_array(4)(190),
      output(5)  => mem_array(5)(190),
      output(6)  => mem_array(6)(190),
      output(7)  => mem_array(7)(190),
      output(8)  => mem_array(8)(190),
      output(9)  => mem_array(9)(190),
      output(10) => mem_array(10)(190),
      output(11) => mem_array(11)(190),
      output(12) => mem_array(12)(190),
      output(13) => mem_array(13)(190),
      output(14) => mem_array(14)(190),
      output(15) => mem_array(15)(190),
      output(16) => mem_array(16)(190),
      output(17) => mem_array(17)(190),
      output(18) => mem_array(18)(190),
      output(19) => mem_array(19)(190),
      output(20) => mem_array(20)(190),
      output(21) => mem_array(21)(190),
      output(22) => mem_array(22)(190),
      output(23) => mem_array(23)(190),
      output(24) => mem_array(24)(190),
      output(25) => mem_array(25)(190),
      output(26) => mem_array(26)(190),
      output(27) => mem_array(27)(190),
      output(28) => mem_array(28)(190),
      output(29) => mem_array(29)(190),
      output(30) => mem_array(30)(190),
      output(31) => mem_array(31)(190),
      output(32) => mem_array(32)(190),
      output(33) => mem_array(33)(190),
      output(34) => mem_array(34)(190),
      output(35) => mem_array(35)(190)
      );
  rom191 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(191),
      output(0)  => mem_array(0)(191),
      output(1)  => mem_array(1)(191),
      output(2)  => mem_array(2)(191),
      output(3)  => mem_array(3)(191),
      output(4)  => mem_array(4)(191),
      output(5)  => mem_array(5)(191),
      output(6)  => mem_array(6)(191),
      output(7)  => mem_array(7)(191),
      output(8)  => mem_array(8)(191),
      output(9)  => mem_array(9)(191),
      output(10) => mem_array(10)(191),
      output(11) => mem_array(11)(191),
      output(12) => mem_array(12)(191),
      output(13) => mem_array(13)(191),
      output(14) => mem_array(14)(191),
      output(15) => mem_array(15)(191),
      output(16) => mem_array(16)(191),
      output(17) => mem_array(17)(191),
      output(18) => mem_array(18)(191),
      output(19) => mem_array(19)(191),
      output(20) => mem_array(20)(191),
      output(21) => mem_array(21)(191),
      output(22) => mem_array(22)(191),
      output(23) => mem_array(23)(191),
      output(24) => mem_array(24)(191),
      output(25) => mem_array(25)(191),
      output(26) => mem_array(26)(191),
      output(27) => mem_array(27)(191),
      output(28) => mem_array(28)(191),
      output(29) => mem_array(29)(191),
      output(30) => mem_array(30)(191),
      output(31) => mem_array(31)(191),
      output(32) => mem_array(32)(191),
      output(33) => mem_array(33)(191),
      output(34) => mem_array(34)(191),
      output(35) => mem_array(35)(191)
      );
  rom192 : entity work.rom
    generic map (
      bits  => 36,
      value => "001011000000000101000000010010100101")
    port map (
      enable_o   => mem_enable_lines(192),
      output(0)  => mem_array(0)(192),
      output(1)  => mem_array(1)(192),
      output(2)  => mem_array(2)(192),
      output(3)  => mem_array(3)(192),
      output(4)  => mem_array(4)(192),
      output(5)  => mem_array(5)(192),
      output(6)  => mem_array(6)(192),
      output(7)  => mem_array(7)(192),
      output(8)  => mem_array(8)(192),
      output(9)  => mem_array(9)(192),
      output(10) => mem_array(10)(192),
      output(11) => mem_array(11)(192),
      output(12) => mem_array(12)(192),
      output(13) => mem_array(13)(192),
      output(14) => mem_array(14)(192),
      output(15) => mem_array(15)(192),
      output(16) => mem_array(16)(192),
      output(17) => mem_array(17)(192),
      output(18) => mem_array(18)(192),
      output(19) => mem_array(19)(192),
      output(20) => mem_array(20)(192),
      output(21) => mem_array(21)(192),
      output(22) => mem_array(22)(192),
      output(23) => mem_array(23)(192),
      output(24) => mem_array(24)(192),
      output(25) => mem_array(25)(192),
      output(26) => mem_array(26)(192),
      output(27) => mem_array(27)(192),
      output(28) => mem_array(28)(192),
      output(29) => mem_array(29)(192),
      output(30) => mem_array(30)(192),
      output(31) => mem_array(31)(192),
      output(32) => mem_array(32)(192),
      output(33) => mem_array(33)(192),
      output(34) => mem_array(34)(192),
      output(35) => mem_array(35)(192)
      );
  rom193 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(193),
      output(0)  => mem_array(0)(193),
      output(1)  => mem_array(1)(193),
      output(2)  => mem_array(2)(193),
      output(3)  => mem_array(3)(193),
      output(4)  => mem_array(4)(193),
      output(5)  => mem_array(5)(193),
      output(6)  => mem_array(6)(193),
      output(7)  => mem_array(7)(193),
      output(8)  => mem_array(8)(193),
      output(9)  => mem_array(9)(193),
      output(10) => mem_array(10)(193),
      output(11) => mem_array(11)(193),
      output(12) => mem_array(12)(193),
      output(13) => mem_array(13)(193),
      output(14) => mem_array(14)(193),
      output(15) => mem_array(15)(193),
      output(16) => mem_array(16)(193),
      output(17) => mem_array(17)(193),
      output(18) => mem_array(18)(193),
      output(19) => mem_array(19)(193),
      output(20) => mem_array(20)(193),
      output(21) => mem_array(21)(193),
      output(22) => mem_array(22)(193),
      output(23) => mem_array(23)(193),
      output(24) => mem_array(24)(193),
      output(25) => mem_array(25)(193),
      output(26) => mem_array(26)(193),
      output(27) => mem_array(27)(193),
      output(28) => mem_array(28)(193),
      output(29) => mem_array(29)(193),
      output(30) => mem_array(30)(193),
      output(31) => mem_array(31)(193),
      output(32) => mem_array(32)(193),
      output(33) => mem_array(33)(193),
      output(34) => mem_array(34)(193),
      output(35) => mem_array(35)(193)
      );
  rom194 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(194),
      output(0)  => mem_array(0)(194),
      output(1)  => mem_array(1)(194),
      output(2)  => mem_array(2)(194),
      output(3)  => mem_array(3)(194),
      output(4)  => mem_array(4)(194),
      output(5)  => mem_array(5)(194),
      output(6)  => mem_array(6)(194),
      output(7)  => mem_array(7)(194),
      output(8)  => mem_array(8)(194),
      output(9)  => mem_array(9)(194),
      output(10) => mem_array(10)(194),
      output(11) => mem_array(11)(194),
      output(12) => mem_array(12)(194),
      output(13) => mem_array(13)(194),
      output(14) => mem_array(14)(194),
      output(15) => mem_array(15)(194),
      output(16) => mem_array(16)(194),
      output(17) => mem_array(17)(194),
      output(18) => mem_array(18)(194),
      output(19) => mem_array(19)(194),
      output(20) => mem_array(20)(194),
      output(21) => mem_array(21)(194),
      output(22) => mem_array(22)(194),
      output(23) => mem_array(23)(194),
      output(24) => mem_array(24)(194),
      output(25) => mem_array(25)(194),
      output(26) => mem_array(26)(194),
      output(27) => mem_array(27)(194),
      output(28) => mem_array(28)(194),
      output(29) => mem_array(29)(194),
      output(30) => mem_array(30)(194),
      output(31) => mem_array(31)(194),
      output(32) => mem_array(32)(194),
      output(33) => mem_array(33)(194),
      output(34) => mem_array(34)(194),
      output(35) => mem_array(35)(194)
      );
  rom195 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(195),
      output(0)  => mem_array(0)(195),
      output(1)  => mem_array(1)(195),
      output(2)  => mem_array(2)(195),
      output(3)  => mem_array(3)(195),
      output(4)  => mem_array(4)(195),
      output(5)  => mem_array(5)(195),
      output(6)  => mem_array(6)(195),
      output(7)  => mem_array(7)(195),
      output(8)  => mem_array(8)(195),
      output(9)  => mem_array(9)(195),
      output(10) => mem_array(10)(195),
      output(11) => mem_array(11)(195),
      output(12) => mem_array(12)(195),
      output(13) => mem_array(13)(195),
      output(14) => mem_array(14)(195),
      output(15) => mem_array(15)(195),
      output(16) => mem_array(16)(195),
      output(17) => mem_array(17)(195),
      output(18) => mem_array(18)(195),
      output(19) => mem_array(19)(195),
      output(20) => mem_array(20)(195),
      output(21) => mem_array(21)(195),
      output(22) => mem_array(22)(195),
      output(23) => mem_array(23)(195),
      output(24) => mem_array(24)(195),
      output(25) => mem_array(25)(195),
      output(26) => mem_array(26)(195),
      output(27) => mem_array(27)(195),
      output(28) => mem_array(28)(195),
      output(29) => mem_array(29)(195),
      output(30) => mem_array(30)(195),
      output(31) => mem_array(31)(195),
      output(32) => mem_array(32)(195),
      output(33) => mem_array(33)(195),
      output(34) => mem_array(34)(195),
      output(35) => mem_array(35)(195)
      );
  rom196 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000100100000110110")
    port map (
      enable_o   => mem_enable_lines(196),
      output(0)  => mem_array(0)(196),
      output(1)  => mem_array(1)(196),
      output(2)  => mem_array(2)(196),
      output(3)  => mem_array(3)(196),
      output(4)  => mem_array(4)(196),
      output(5)  => mem_array(5)(196),
      output(6)  => mem_array(6)(196),
      output(7)  => mem_array(7)(196),
      output(8)  => mem_array(8)(196),
      output(9)  => mem_array(9)(196),
      output(10) => mem_array(10)(196),
      output(11) => mem_array(11)(196),
      output(12) => mem_array(12)(196),
      output(13) => mem_array(13)(196),
      output(14) => mem_array(14)(196),
      output(15) => mem_array(15)(196),
      output(16) => mem_array(16)(196),
      output(17) => mem_array(17)(196),
      output(18) => mem_array(18)(196),
      output(19) => mem_array(19)(196),
      output(20) => mem_array(20)(196),
      output(21) => mem_array(21)(196),
      output(22) => mem_array(22)(196),
      output(23) => mem_array(23)(196),
      output(24) => mem_array(24)(196),
      output(25) => mem_array(25)(196),
      output(26) => mem_array(26)(196),
      output(27) => mem_array(27)(196),
      output(28) => mem_array(28)(196),
      output(29) => mem_array(29)(196),
      output(30) => mem_array(30)(196),
      output(31) => mem_array(31)(196),
      output(32) => mem_array(32)(196),
      output(33) => mem_array(33)(196),
      output(34) => mem_array(34)(196),
      output(35) => mem_array(35)(196)
      );
  rom197 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001001010010000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(197),
      output(0)  => mem_array(0)(197),
      output(1)  => mem_array(1)(197),
      output(2)  => mem_array(2)(197),
      output(3)  => mem_array(3)(197),
      output(4)  => mem_array(4)(197),
      output(5)  => mem_array(5)(197),
      output(6)  => mem_array(6)(197),
      output(7)  => mem_array(7)(197),
      output(8)  => mem_array(8)(197),
      output(9)  => mem_array(9)(197),
      output(10) => mem_array(10)(197),
      output(11) => mem_array(11)(197),
      output(12) => mem_array(12)(197),
      output(13) => mem_array(13)(197),
      output(14) => mem_array(14)(197),
      output(15) => mem_array(15)(197),
      output(16) => mem_array(16)(197),
      output(17) => mem_array(17)(197),
      output(18) => mem_array(18)(197),
      output(19) => mem_array(19)(197),
      output(20) => mem_array(20)(197),
      output(21) => mem_array(21)(197),
      output(22) => mem_array(22)(197),
      output(23) => mem_array(23)(197),
      output(24) => mem_array(24)(197),
      output(25) => mem_array(25)(197),
      output(26) => mem_array(26)(197),
      output(27) => mem_array(27)(197),
      output(28) => mem_array(28)(197),
      output(29) => mem_array(29)(197),
      output(30) => mem_array(30)(197),
      output(31) => mem_array(31)(197),
      output(32) => mem_array(32)(197),
      output(33) => mem_array(33)(197),
      output(34) => mem_array(34)(197),
      output(35) => mem_array(35)(197)
      );
  rom198 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(198),
      output(0)  => mem_array(0)(198),
      output(1)  => mem_array(1)(198),
      output(2)  => mem_array(2)(198),
      output(3)  => mem_array(3)(198),
      output(4)  => mem_array(4)(198),
      output(5)  => mem_array(5)(198),
      output(6)  => mem_array(6)(198),
      output(7)  => mem_array(7)(198),
      output(8)  => mem_array(8)(198),
      output(9)  => mem_array(9)(198),
      output(10) => mem_array(10)(198),
      output(11) => mem_array(11)(198),
      output(12) => mem_array(12)(198),
      output(13) => mem_array(13)(198),
      output(14) => mem_array(14)(198),
      output(15) => mem_array(15)(198),
      output(16) => mem_array(16)(198),
      output(17) => mem_array(17)(198),
      output(18) => mem_array(18)(198),
      output(19) => mem_array(19)(198),
      output(20) => mem_array(20)(198),
      output(21) => mem_array(21)(198),
      output(22) => mem_array(22)(198),
      output(23) => mem_array(23)(198),
      output(24) => mem_array(24)(198),
      output(25) => mem_array(25)(198),
      output(26) => mem_array(26)(198),
      output(27) => mem_array(27)(198),
      output(28) => mem_array(28)(198),
      output(29) => mem_array(29)(198),
      output(30) => mem_array(30)(198),
      output(31) => mem_array(31)(198),
      output(32) => mem_array(32)(198),
      output(33) => mem_array(33)(198),
      output(34) => mem_array(34)(198),
      output(35) => mem_array(35)(198)
      );
  rom199 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(199),
      output(0)  => mem_array(0)(199),
      output(1)  => mem_array(1)(199),
      output(2)  => mem_array(2)(199),
      output(3)  => mem_array(3)(199),
      output(4)  => mem_array(4)(199),
      output(5)  => mem_array(5)(199),
      output(6)  => mem_array(6)(199),
      output(7)  => mem_array(7)(199),
      output(8)  => mem_array(8)(199),
      output(9)  => mem_array(9)(199),
      output(10) => mem_array(10)(199),
      output(11) => mem_array(11)(199),
      output(12) => mem_array(12)(199),
      output(13) => mem_array(13)(199),
      output(14) => mem_array(14)(199),
      output(15) => mem_array(15)(199),
      output(16) => mem_array(16)(199),
      output(17) => mem_array(17)(199),
      output(18) => mem_array(18)(199),
      output(19) => mem_array(19)(199),
      output(20) => mem_array(20)(199),
      output(21) => mem_array(21)(199),
      output(22) => mem_array(22)(199),
      output(23) => mem_array(23)(199),
      output(24) => mem_array(24)(199),
      output(25) => mem_array(25)(199),
      output(26) => mem_array(26)(199),
      output(27) => mem_array(27)(199),
      output(28) => mem_array(28)(199),
      output(29) => mem_array(29)(199),
      output(30) => mem_array(30)(199),
      output(31) => mem_array(31)(199),
      output(32) => mem_array(32)(199),
      output(33) => mem_array(33)(199),
      output(34) => mem_array(34)(199),
      output(35) => mem_array(35)(199)
      );
  rom200 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(200),
      output(0)  => mem_array(0)(200),
      output(1)  => mem_array(1)(200),
      output(2)  => mem_array(2)(200),
      output(3)  => mem_array(3)(200),
      output(4)  => mem_array(4)(200),
      output(5)  => mem_array(5)(200),
      output(6)  => mem_array(6)(200),
      output(7)  => mem_array(7)(200),
      output(8)  => mem_array(8)(200),
      output(9)  => mem_array(9)(200),
      output(10) => mem_array(10)(200),
      output(11) => mem_array(11)(200),
      output(12) => mem_array(12)(200),
      output(13) => mem_array(13)(200),
      output(14) => mem_array(14)(200),
      output(15) => mem_array(15)(200),
      output(16) => mem_array(16)(200),
      output(17) => mem_array(17)(200),
      output(18) => mem_array(18)(200),
      output(19) => mem_array(19)(200),
      output(20) => mem_array(20)(200),
      output(21) => mem_array(21)(200),
      output(22) => mem_array(22)(200),
      output(23) => mem_array(23)(200),
      output(24) => mem_array(24)(200),
      output(25) => mem_array(25)(200),
      output(26) => mem_array(26)(200),
      output(27) => mem_array(27)(200),
      output(28) => mem_array(28)(200),
      output(29) => mem_array(29)(200),
      output(30) => mem_array(30)(200),
      output(31) => mem_array(31)(200),
      output(32) => mem_array(32)(200),
      output(33) => mem_array(33)(200),
      output(34) => mem_array(34)(200),
      output(35) => mem_array(35)(200)
      );
  rom201 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(201),
      output(0)  => mem_array(0)(201),
      output(1)  => mem_array(1)(201),
      output(2)  => mem_array(2)(201),
      output(3)  => mem_array(3)(201),
      output(4)  => mem_array(4)(201),
      output(5)  => mem_array(5)(201),
      output(6)  => mem_array(6)(201),
      output(7)  => mem_array(7)(201),
      output(8)  => mem_array(8)(201),
      output(9)  => mem_array(9)(201),
      output(10) => mem_array(10)(201),
      output(11) => mem_array(11)(201),
      output(12) => mem_array(12)(201),
      output(13) => mem_array(13)(201),
      output(14) => mem_array(14)(201),
      output(15) => mem_array(15)(201),
      output(16) => mem_array(16)(201),
      output(17) => mem_array(17)(201),
      output(18) => mem_array(18)(201),
      output(19) => mem_array(19)(201),
      output(20) => mem_array(20)(201),
      output(21) => mem_array(21)(201),
      output(22) => mem_array(22)(201),
      output(23) => mem_array(23)(201),
      output(24) => mem_array(24)(201),
      output(25) => mem_array(25)(201),
      output(26) => mem_array(26)(201),
      output(27) => mem_array(27)(201),
      output(28) => mem_array(28)(201),
      output(29) => mem_array(29)(201),
      output(30) => mem_array(30)(201),
      output(31) => mem_array(31)(201),
      output(32) => mem_array(32)(201),
      output(33) => mem_array(33)(201),
      output(34) => mem_array(34)(201),
      output(35) => mem_array(35)(201)
      );
  rom202 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(202),
      output(0)  => mem_array(0)(202),
      output(1)  => mem_array(1)(202),
      output(2)  => mem_array(2)(202),
      output(3)  => mem_array(3)(202),
      output(4)  => mem_array(4)(202),
      output(5)  => mem_array(5)(202),
      output(6)  => mem_array(6)(202),
      output(7)  => mem_array(7)(202),
      output(8)  => mem_array(8)(202),
      output(9)  => mem_array(9)(202),
      output(10) => mem_array(10)(202),
      output(11) => mem_array(11)(202),
      output(12) => mem_array(12)(202),
      output(13) => mem_array(13)(202),
      output(14) => mem_array(14)(202),
      output(15) => mem_array(15)(202),
      output(16) => mem_array(16)(202),
      output(17) => mem_array(17)(202),
      output(18) => mem_array(18)(202),
      output(19) => mem_array(19)(202),
      output(20) => mem_array(20)(202),
      output(21) => mem_array(21)(202),
      output(22) => mem_array(22)(202),
      output(23) => mem_array(23)(202),
      output(24) => mem_array(24)(202),
      output(25) => mem_array(25)(202),
      output(26) => mem_array(26)(202),
      output(27) => mem_array(27)(202),
      output(28) => mem_array(28)(202),
      output(29) => mem_array(29)(202),
      output(30) => mem_array(30)(202),
      output(31) => mem_array(31)(202),
      output(32) => mem_array(32)(202),
      output(33) => mem_array(33)(202),
      output(34) => mem_array(34)(202),
      output(35) => mem_array(35)(202)
      );
  rom203 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000100001000000110101000000100001")
    port map (
      enable_o   => mem_enable_lines(203),
      output(0)  => mem_array(0)(203),
      output(1)  => mem_array(1)(203),
      output(2)  => mem_array(2)(203),
      output(3)  => mem_array(3)(203),
      output(4)  => mem_array(4)(203),
      output(5)  => mem_array(5)(203),
      output(6)  => mem_array(6)(203),
      output(7)  => mem_array(7)(203),
      output(8)  => mem_array(8)(203),
      output(9)  => mem_array(9)(203),
      output(10) => mem_array(10)(203),
      output(11) => mem_array(11)(203),
      output(12) => mem_array(12)(203),
      output(13) => mem_array(13)(203),
      output(14) => mem_array(14)(203),
      output(15) => mem_array(15)(203),
      output(16) => mem_array(16)(203),
      output(17) => mem_array(17)(203),
      output(18) => mem_array(18)(203),
      output(19) => mem_array(19)(203),
      output(20) => mem_array(20)(203),
      output(21) => mem_array(21)(203),
      output(22) => mem_array(22)(203),
      output(23) => mem_array(23)(203),
      output(24) => mem_array(24)(203),
      output(25) => mem_array(25)(203),
      output(26) => mem_array(26)(203),
      output(27) => mem_array(27)(203),
      output(28) => mem_array(28)(203),
      output(29) => mem_array(29)(203),
      output(30) => mem_array(30)(203),
      output(31) => mem_array(31)(203),
      output(32) => mem_array(32)(203),
      output(33) => mem_array(33)(203),
      output(34) => mem_array(34)(203),
      output(35) => mem_array(35)(203)
      );
  rom204 : entity work.rom
    generic map (
      bits  => 36,
      value => "000100000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(204),
      output(0)  => mem_array(0)(204),
      output(1)  => mem_array(1)(204),
      output(2)  => mem_array(2)(204),
      output(3)  => mem_array(3)(204),
      output(4)  => mem_array(4)(204),
      output(5)  => mem_array(5)(204),
      output(6)  => mem_array(6)(204),
      output(7)  => mem_array(7)(204),
      output(8)  => mem_array(8)(204),
      output(9)  => mem_array(9)(204),
      output(10) => mem_array(10)(204),
      output(11) => mem_array(11)(204),
      output(12) => mem_array(12)(204),
      output(13) => mem_array(13)(204),
      output(14) => mem_array(14)(204),
      output(15) => mem_array(15)(204),
      output(16) => mem_array(16)(204),
      output(17) => mem_array(17)(204),
      output(18) => mem_array(18)(204),
      output(19) => mem_array(19)(204),
      output(20) => mem_array(20)(204),
      output(21) => mem_array(21)(204),
      output(22) => mem_array(22)(204),
      output(23) => mem_array(23)(204),
      output(24) => mem_array(24)(204),
      output(25) => mem_array(25)(204),
      output(26) => mem_array(26)(204),
      output(27) => mem_array(27)(204),
      output(28) => mem_array(28)(204),
      output(29) => mem_array(29)(204),
      output(30) => mem_array(30)(204),
      output(31) => mem_array(31)(204),
      output(32) => mem_array(32)(204),
      output(33) => mem_array(33)(204),
      output(34) => mem_array(34)(204),
      output(35) => mem_array(35)(204)
      );
  rom205 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(205),
      output(0)  => mem_array(0)(205),
      output(1)  => mem_array(1)(205),
      output(2)  => mem_array(2)(205),
      output(3)  => mem_array(3)(205),
      output(4)  => mem_array(4)(205),
      output(5)  => mem_array(5)(205),
      output(6)  => mem_array(6)(205),
      output(7)  => mem_array(7)(205),
      output(8)  => mem_array(8)(205),
      output(9)  => mem_array(9)(205),
      output(10) => mem_array(10)(205),
      output(11) => mem_array(11)(205),
      output(12) => mem_array(12)(205),
      output(13) => mem_array(13)(205),
      output(14) => mem_array(14)(205),
      output(15) => mem_array(15)(205),
      output(16) => mem_array(16)(205),
      output(17) => mem_array(17)(205),
      output(18) => mem_array(18)(205),
      output(19) => mem_array(19)(205),
      output(20) => mem_array(20)(205),
      output(21) => mem_array(21)(205),
      output(22) => mem_array(22)(205),
      output(23) => mem_array(23)(205),
      output(24) => mem_array(24)(205),
      output(25) => mem_array(25)(205),
      output(26) => mem_array(26)(205),
      output(27) => mem_array(27)(205),
      output(28) => mem_array(28)(205),
      output(29) => mem_array(29)(205),
      output(30) => mem_array(30)(205),
      output(31) => mem_array(31)(205),
      output(32) => mem_array(32)(205),
      output(33) => mem_array(33)(205),
      output(34) => mem_array(34)(205),
      output(35) => mem_array(35)(205)
      );
  rom206 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(206),
      output(0)  => mem_array(0)(206),
      output(1)  => mem_array(1)(206),
      output(2)  => mem_array(2)(206),
      output(3)  => mem_array(3)(206),
      output(4)  => mem_array(4)(206),
      output(5)  => mem_array(5)(206),
      output(6)  => mem_array(6)(206),
      output(7)  => mem_array(7)(206),
      output(8)  => mem_array(8)(206),
      output(9)  => mem_array(9)(206),
      output(10) => mem_array(10)(206),
      output(11) => mem_array(11)(206),
      output(12) => mem_array(12)(206),
      output(13) => mem_array(13)(206),
      output(14) => mem_array(14)(206),
      output(15) => mem_array(15)(206),
      output(16) => mem_array(16)(206),
      output(17) => mem_array(17)(206),
      output(18) => mem_array(18)(206),
      output(19) => mem_array(19)(206),
      output(20) => mem_array(20)(206),
      output(21) => mem_array(21)(206),
      output(22) => mem_array(22)(206),
      output(23) => mem_array(23)(206),
      output(24) => mem_array(24)(206),
      output(25) => mem_array(25)(206),
      output(26) => mem_array(26)(206),
      output(27) => mem_array(27)(206),
      output(28) => mem_array(28)(206),
      output(29) => mem_array(29)(206),
      output(30) => mem_array(30)(206),
      output(31) => mem_array(31)(206),
      output(32) => mem_array(32)(206),
      output(33) => mem_array(33)(206),
      output(34) => mem_array(34)(206),
      output(35) => mem_array(35)(206)
      );
  rom207 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(207),
      output(0)  => mem_array(0)(207),
      output(1)  => mem_array(1)(207),
      output(2)  => mem_array(2)(207),
      output(3)  => mem_array(3)(207),
      output(4)  => mem_array(4)(207),
      output(5)  => mem_array(5)(207),
      output(6)  => mem_array(6)(207),
      output(7)  => mem_array(7)(207),
      output(8)  => mem_array(8)(207),
      output(9)  => mem_array(9)(207),
      output(10) => mem_array(10)(207),
      output(11) => mem_array(11)(207),
      output(12) => mem_array(12)(207),
      output(13) => mem_array(13)(207),
      output(14) => mem_array(14)(207),
      output(15) => mem_array(15)(207),
      output(16) => mem_array(16)(207),
      output(17) => mem_array(17)(207),
      output(18) => mem_array(18)(207),
      output(19) => mem_array(19)(207),
      output(20) => mem_array(20)(207),
      output(21) => mem_array(21)(207),
      output(22) => mem_array(22)(207),
      output(23) => mem_array(23)(207),
      output(24) => mem_array(24)(207),
      output(25) => mem_array(25)(207),
      output(26) => mem_array(26)(207),
      output(27) => mem_array(27)(207),
      output(28) => mem_array(28)(207),
      output(29) => mem_array(29)(207),
      output(30) => mem_array(30)(207),
      output(31) => mem_array(31)(207),
      output(32) => mem_array(32)(207),
      output(33) => mem_array(33)(207),
      output(34) => mem_array(34)(207),
      output(35) => mem_array(35)(207)
      );
  rom208 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(208),
      output(0)  => mem_array(0)(208),
      output(1)  => mem_array(1)(208),
      output(2)  => mem_array(2)(208),
      output(3)  => mem_array(3)(208),
      output(4)  => mem_array(4)(208),
      output(5)  => mem_array(5)(208),
      output(6)  => mem_array(6)(208),
      output(7)  => mem_array(7)(208),
      output(8)  => mem_array(8)(208),
      output(9)  => mem_array(9)(208),
      output(10) => mem_array(10)(208),
      output(11) => mem_array(11)(208),
      output(12) => mem_array(12)(208),
      output(13) => mem_array(13)(208),
      output(14) => mem_array(14)(208),
      output(15) => mem_array(15)(208),
      output(16) => mem_array(16)(208),
      output(17) => mem_array(17)(208),
      output(18) => mem_array(18)(208),
      output(19) => mem_array(19)(208),
      output(20) => mem_array(20)(208),
      output(21) => mem_array(21)(208),
      output(22) => mem_array(22)(208),
      output(23) => mem_array(23)(208),
      output(24) => mem_array(24)(208),
      output(25) => mem_array(25)(208),
      output(26) => mem_array(26)(208),
      output(27) => mem_array(27)(208),
      output(28) => mem_array(28)(208),
      output(29) => mem_array(29)(208),
      output(30) => mem_array(30)(208),
      output(31) => mem_array(31)(208),
      output(32) => mem_array(32)(208),
      output(33) => mem_array(33)(208),
      output(34) => mem_array(34)(208),
      output(35) => mem_array(35)(208)
      );
  rom209 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(209),
      output(0)  => mem_array(0)(209),
      output(1)  => mem_array(1)(209),
      output(2)  => mem_array(2)(209),
      output(3)  => mem_array(3)(209),
      output(4)  => mem_array(4)(209),
      output(5)  => mem_array(5)(209),
      output(6)  => mem_array(6)(209),
      output(7)  => mem_array(7)(209),
      output(8)  => mem_array(8)(209),
      output(9)  => mem_array(9)(209),
      output(10) => mem_array(10)(209),
      output(11) => mem_array(11)(209),
      output(12) => mem_array(12)(209),
      output(13) => mem_array(13)(209),
      output(14) => mem_array(14)(209),
      output(15) => mem_array(15)(209),
      output(16) => mem_array(16)(209),
      output(17) => mem_array(17)(209),
      output(18) => mem_array(18)(209),
      output(19) => mem_array(19)(209),
      output(20) => mem_array(20)(209),
      output(21) => mem_array(21)(209),
      output(22) => mem_array(22)(209),
      output(23) => mem_array(23)(209),
      output(24) => mem_array(24)(209),
      output(25) => mem_array(25)(209),
      output(26) => mem_array(26)(209),
      output(27) => mem_array(27)(209),
      output(28) => mem_array(28)(209),
      output(29) => mem_array(29)(209),
      output(30) => mem_array(30)(209),
      output(31) => mem_array(31)(209),
      output(32) => mem_array(32)(209),
      output(33) => mem_array(33)(209),
      output(34) => mem_array(34)(209),
      output(35) => mem_array(35)(209)
      );
  rom210 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(210),
      output(0)  => mem_array(0)(210),
      output(1)  => mem_array(1)(210),
      output(2)  => mem_array(2)(210),
      output(3)  => mem_array(3)(210),
      output(4)  => mem_array(4)(210),
      output(5)  => mem_array(5)(210),
      output(6)  => mem_array(6)(210),
      output(7)  => mem_array(7)(210),
      output(8)  => mem_array(8)(210),
      output(9)  => mem_array(9)(210),
      output(10) => mem_array(10)(210),
      output(11) => mem_array(11)(210),
      output(12) => mem_array(12)(210),
      output(13) => mem_array(13)(210),
      output(14) => mem_array(14)(210),
      output(15) => mem_array(15)(210),
      output(16) => mem_array(16)(210),
      output(17) => mem_array(17)(210),
      output(18) => mem_array(18)(210),
      output(19) => mem_array(19)(210),
      output(20) => mem_array(20)(210),
      output(21) => mem_array(21)(210),
      output(22) => mem_array(22)(210),
      output(23) => mem_array(23)(210),
      output(24) => mem_array(24)(210),
      output(25) => mem_array(25)(210),
      output(26) => mem_array(26)(210),
      output(27) => mem_array(27)(210),
      output(28) => mem_array(28)(210),
      output(29) => mem_array(29)(210),
      output(30) => mem_array(30)(210),
      output(31) => mem_array(31)(210),
      output(32) => mem_array(32)(210),
      output(33) => mem_array(33)(210),
      output(34) => mem_array(34)(210),
      output(35) => mem_array(35)(210)
      );
  rom211 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(211),
      output(0)  => mem_array(0)(211),
      output(1)  => mem_array(1)(211),
      output(2)  => mem_array(2)(211),
      output(3)  => mem_array(3)(211),
      output(4)  => mem_array(4)(211),
      output(5)  => mem_array(5)(211),
      output(6)  => mem_array(6)(211),
      output(7)  => mem_array(7)(211),
      output(8)  => mem_array(8)(211),
      output(9)  => mem_array(9)(211),
      output(10) => mem_array(10)(211),
      output(11) => mem_array(11)(211),
      output(12) => mem_array(12)(211),
      output(13) => mem_array(13)(211),
      output(14) => mem_array(14)(211),
      output(15) => mem_array(15)(211),
      output(16) => mem_array(16)(211),
      output(17) => mem_array(17)(211),
      output(18) => mem_array(18)(211),
      output(19) => mem_array(19)(211),
      output(20) => mem_array(20)(211),
      output(21) => mem_array(21)(211),
      output(22) => mem_array(22)(211),
      output(23) => mem_array(23)(211),
      output(24) => mem_array(24)(211),
      output(25) => mem_array(25)(211),
      output(26) => mem_array(26)(211),
      output(27) => mem_array(27)(211),
      output(28) => mem_array(28)(211),
      output(29) => mem_array(29)(211),
      output(30) => mem_array(30)(211),
      output(31) => mem_array(31)(211),
      output(32) => mem_array(32)(211),
      output(33) => mem_array(33)(211),
      output(34) => mem_array(34)(211),
      output(35) => mem_array(35)(211)
      );
  rom212 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(212),
      output(0)  => mem_array(0)(212),
      output(1)  => mem_array(1)(212),
      output(2)  => mem_array(2)(212),
      output(3)  => mem_array(3)(212),
      output(4)  => mem_array(4)(212),
      output(5)  => mem_array(5)(212),
      output(6)  => mem_array(6)(212),
      output(7)  => mem_array(7)(212),
      output(8)  => mem_array(8)(212),
      output(9)  => mem_array(9)(212),
      output(10) => mem_array(10)(212),
      output(11) => mem_array(11)(212),
      output(12) => mem_array(12)(212),
      output(13) => mem_array(13)(212),
      output(14) => mem_array(14)(212),
      output(15) => mem_array(15)(212),
      output(16) => mem_array(16)(212),
      output(17) => mem_array(17)(212),
      output(18) => mem_array(18)(212),
      output(19) => mem_array(19)(212),
      output(20) => mem_array(20)(212),
      output(21) => mem_array(21)(212),
      output(22) => mem_array(22)(212),
      output(23) => mem_array(23)(212),
      output(24) => mem_array(24)(212),
      output(25) => mem_array(25)(212),
      output(26) => mem_array(26)(212),
      output(27) => mem_array(27)(212),
      output(28) => mem_array(28)(212),
      output(29) => mem_array(29)(212),
      output(30) => mem_array(30)(212),
      output(31) => mem_array(31)(212),
      output(32) => mem_array(32)(212),
      output(33) => mem_array(33)(212),
      output(34) => mem_array(34)(212),
      output(35) => mem_array(35)(212)
      );
  rom213 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(213),
      output(0)  => mem_array(0)(213),
      output(1)  => mem_array(1)(213),
      output(2)  => mem_array(2)(213),
      output(3)  => mem_array(3)(213),
      output(4)  => mem_array(4)(213),
      output(5)  => mem_array(5)(213),
      output(6)  => mem_array(6)(213),
      output(7)  => mem_array(7)(213),
      output(8)  => mem_array(8)(213),
      output(9)  => mem_array(9)(213),
      output(10) => mem_array(10)(213),
      output(11) => mem_array(11)(213),
      output(12) => mem_array(12)(213),
      output(13) => mem_array(13)(213),
      output(14) => mem_array(14)(213),
      output(15) => mem_array(15)(213),
      output(16) => mem_array(16)(213),
      output(17) => mem_array(17)(213),
      output(18) => mem_array(18)(213),
      output(19) => mem_array(19)(213),
      output(20) => mem_array(20)(213),
      output(21) => mem_array(21)(213),
      output(22) => mem_array(22)(213),
      output(23) => mem_array(23)(213),
      output(24) => mem_array(24)(213),
      output(25) => mem_array(25)(213),
      output(26) => mem_array(26)(213),
      output(27) => mem_array(27)(213),
      output(28) => mem_array(28)(213),
      output(29) => mem_array(29)(213),
      output(30) => mem_array(30)(213),
      output(31) => mem_array(31)(213),
      output(32) => mem_array(32)(213),
      output(33) => mem_array(33)(213),
      output(34) => mem_array(34)(213),
      output(35) => mem_array(35)(213)
      );
  rom214 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(214),
      output(0)  => mem_array(0)(214),
      output(1)  => mem_array(1)(214),
      output(2)  => mem_array(2)(214),
      output(3)  => mem_array(3)(214),
      output(4)  => mem_array(4)(214),
      output(5)  => mem_array(5)(214),
      output(6)  => mem_array(6)(214),
      output(7)  => mem_array(7)(214),
      output(8)  => mem_array(8)(214),
      output(9)  => mem_array(9)(214),
      output(10) => mem_array(10)(214),
      output(11) => mem_array(11)(214),
      output(12) => mem_array(12)(214),
      output(13) => mem_array(13)(214),
      output(14) => mem_array(14)(214),
      output(15) => mem_array(15)(214),
      output(16) => mem_array(16)(214),
      output(17) => mem_array(17)(214),
      output(18) => mem_array(18)(214),
      output(19) => mem_array(19)(214),
      output(20) => mem_array(20)(214),
      output(21) => mem_array(21)(214),
      output(22) => mem_array(22)(214),
      output(23) => mem_array(23)(214),
      output(24) => mem_array(24)(214),
      output(25) => mem_array(25)(214),
      output(26) => mem_array(26)(214),
      output(27) => mem_array(27)(214),
      output(28) => mem_array(28)(214),
      output(29) => mem_array(29)(214),
      output(30) => mem_array(30)(214),
      output(31) => mem_array(31)(214),
      output(32) => mem_array(32)(214),
      output(33) => mem_array(33)(214),
      output(34) => mem_array(34)(214),
      output(35) => mem_array(35)(214)
      );
  rom215 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(215),
      output(0)  => mem_array(0)(215),
      output(1)  => mem_array(1)(215),
      output(2)  => mem_array(2)(215),
      output(3)  => mem_array(3)(215),
      output(4)  => mem_array(4)(215),
      output(5)  => mem_array(5)(215),
      output(6)  => mem_array(6)(215),
      output(7)  => mem_array(7)(215),
      output(8)  => mem_array(8)(215),
      output(9)  => mem_array(9)(215),
      output(10) => mem_array(10)(215),
      output(11) => mem_array(11)(215),
      output(12) => mem_array(12)(215),
      output(13) => mem_array(13)(215),
      output(14) => mem_array(14)(215),
      output(15) => mem_array(15)(215),
      output(16) => mem_array(16)(215),
      output(17) => mem_array(17)(215),
      output(18) => mem_array(18)(215),
      output(19) => mem_array(19)(215),
      output(20) => mem_array(20)(215),
      output(21) => mem_array(21)(215),
      output(22) => mem_array(22)(215),
      output(23) => mem_array(23)(215),
      output(24) => mem_array(24)(215),
      output(25) => mem_array(25)(215),
      output(26) => mem_array(26)(215),
      output(27) => mem_array(27)(215),
      output(28) => mem_array(28)(215),
      output(29) => mem_array(29)(215),
      output(30) => mem_array(30)(215),
      output(31) => mem_array(31)(215),
      output(32) => mem_array(32)(215),
      output(33) => mem_array(33)(215),
      output(34) => mem_array(34)(215),
      output(35) => mem_array(35)(215)
      );
  rom216 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(216),
      output(0)  => mem_array(0)(216),
      output(1)  => mem_array(1)(216),
      output(2)  => mem_array(2)(216),
      output(3)  => mem_array(3)(216),
      output(4)  => mem_array(4)(216),
      output(5)  => mem_array(5)(216),
      output(6)  => mem_array(6)(216),
      output(7)  => mem_array(7)(216),
      output(8)  => mem_array(8)(216),
      output(9)  => mem_array(9)(216),
      output(10) => mem_array(10)(216),
      output(11) => mem_array(11)(216),
      output(12) => mem_array(12)(216),
      output(13) => mem_array(13)(216),
      output(14) => mem_array(14)(216),
      output(15) => mem_array(15)(216),
      output(16) => mem_array(16)(216),
      output(17) => mem_array(17)(216),
      output(18) => mem_array(18)(216),
      output(19) => mem_array(19)(216),
      output(20) => mem_array(20)(216),
      output(21) => mem_array(21)(216),
      output(22) => mem_array(22)(216),
      output(23) => mem_array(23)(216),
      output(24) => mem_array(24)(216),
      output(25) => mem_array(25)(216),
      output(26) => mem_array(26)(216),
      output(27) => mem_array(27)(216),
      output(28) => mem_array(28)(216),
      output(29) => mem_array(29)(216),
      output(30) => mem_array(30)(216),
      output(31) => mem_array(31)(216),
      output(32) => mem_array(32)(216),
      output(33) => mem_array(33)(216),
      output(34) => mem_array(34)(216),
      output(35) => mem_array(35)(216)
      );
  rom217 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(217),
      output(0)  => mem_array(0)(217),
      output(1)  => mem_array(1)(217),
      output(2)  => mem_array(2)(217),
      output(3)  => mem_array(3)(217),
      output(4)  => mem_array(4)(217),
      output(5)  => mem_array(5)(217),
      output(6)  => mem_array(6)(217),
      output(7)  => mem_array(7)(217),
      output(8)  => mem_array(8)(217),
      output(9)  => mem_array(9)(217),
      output(10) => mem_array(10)(217),
      output(11) => mem_array(11)(217),
      output(12) => mem_array(12)(217),
      output(13) => mem_array(13)(217),
      output(14) => mem_array(14)(217),
      output(15) => mem_array(15)(217),
      output(16) => mem_array(16)(217),
      output(17) => mem_array(17)(217),
      output(18) => mem_array(18)(217),
      output(19) => mem_array(19)(217),
      output(20) => mem_array(20)(217),
      output(21) => mem_array(21)(217),
      output(22) => mem_array(22)(217),
      output(23) => mem_array(23)(217),
      output(24) => mem_array(24)(217),
      output(25) => mem_array(25)(217),
      output(26) => mem_array(26)(217),
      output(27) => mem_array(27)(217),
      output(28) => mem_array(28)(217),
      output(29) => mem_array(29)(217),
      output(30) => mem_array(30)(217),
      output(31) => mem_array(31)(217),
      output(32) => mem_array(32)(217),
      output(33) => mem_array(33)(217),
      output(34) => mem_array(34)(217),
      output(35) => mem_array(35)(217)
      );
  rom218 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000100000000100")
    port map (
      enable_o   => mem_enable_lines(218),
      output(0)  => mem_array(0)(218),
      output(1)  => mem_array(1)(218),
      output(2)  => mem_array(2)(218),
      output(3)  => mem_array(3)(218),
      output(4)  => mem_array(4)(218),
      output(5)  => mem_array(5)(218),
      output(6)  => mem_array(6)(218),
      output(7)  => mem_array(7)(218),
      output(8)  => mem_array(8)(218),
      output(9)  => mem_array(9)(218),
      output(10) => mem_array(10)(218),
      output(11) => mem_array(11)(218),
      output(12) => mem_array(12)(218),
      output(13) => mem_array(13)(218),
      output(14) => mem_array(14)(218),
      output(15) => mem_array(15)(218),
      output(16) => mem_array(16)(218),
      output(17) => mem_array(17)(218),
      output(18) => mem_array(18)(218),
      output(19) => mem_array(19)(218),
      output(20) => mem_array(20)(218),
      output(21) => mem_array(21)(218),
      output(22) => mem_array(22)(218),
      output(23) => mem_array(23)(218),
      output(24) => mem_array(24)(218),
      output(25) => mem_array(25)(218),
      output(26) => mem_array(26)(218),
      output(27) => mem_array(27)(218),
      output(28) => mem_array(28)(218),
      output(29) => mem_array(29)(218),
      output(30) => mem_array(30)(218),
      output(31) => mem_array(31)(218),
      output(32) => mem_array(32)(218),
      output(33) => mem_array(33)(218),
      output(34) => mem_array(34)(218),
      output(35) => mem_array(35)(218)
      );
  rom219 : entity work.rom
    generic map (
      bits  => 36,
      value => "001101010000001000010001000001111111")
    port map (
      enable_o   => mem_enable_lines(219),
      output(0)  => mem_array(0)(219),
      output(1)  => mem_array(1)(219),
      output(2)  => mem_array(2)(219),
      output(3)  => mem_array(3)(219),
      output(4)  => mem_array(4)(219),
      output(5)  => mem_array(5)(219),
      output(6)  => mem_array(6)(219),
      output(7)  => mem_array(7)(219),
      output(8)  => mem_array(8)(219),
      output(9)  => mem_array(9)(219),
      output(10) => mem_array(10)(219),
      output(11) => mem_array(11)(219),
      output(12) => mem_array(12)(219),
      output(13) => mem_array(13)(219),
      output(14) => mem_array(14)(219),
      output(15) => mem_array(15)(219),
      output(16) => mem_array(16)(219),
      output(17) => mem_array(17)(219),
      output(18) => mem_array(18)(219),
      output(19) => mem_array(19)(219),
      output(20) => mem_array(20)(219),
      output(21) => mem_array(21)(219),
      output(22) => mem_array(22)(219),
      output(23) => mem_array(23)(219),
      output(24) => mem_array(24)(219),
      output(25) => mem_array(25)(219),
      output(26) => mem_array(26)(219),
      output(27) => mem_array(27)(219),
      output(28) => mem_array(28)(219),
      output(29) => mem_array(29)(219),
      output(30) => mem_array(30)(219),
      output(31) => mem_array(31)(219),
      output(32) => mem_array(32)(219),
      output(33) => mem_array(33)(219),
      output(34) => mem_array(34)(219),
      output(35) => mem_array(35)(219)
      );
  rom220 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(220),
      output(0)  => mem_array(0)(220),
      output(1)  => mem_array(1)(220),
      output(2)  => mem_array(2)(220),
      output(3)  => mem_array(3)(220),
      output(4)  => mem_array(4)(220),
      output(5)  => mem_array(5)(220),
      output(6)  => mem_array(6)(220),
      output(7)  => mem_array(7)(220),
      output(8)  => mem_array(8)(220),
      output(9)  => mem_array(9)(220),
      output(10) => mem_array(10)(220),
      output(11) => mem_array(11)(220),
      output(12) => mem_array(12)(220),
      output(13) => mem_array(13)(220),
      output(14) => mem_array(14)(220),
      output(15) => mem_array(15)(220),
      output(16) => mem_array(16)(220),
      output(17) => mem_array(17)(220),
      output(18) => mem_array(18)(220),
      output(19) => mem_array(19)(220),
      output(20) => mem_array(20)(220),
      output(21) => mem_array(21)(220),
      output(22) => mem_array(22)(220),
      output(23) => mem_array(23)(220),
      output(24) => mem_array(24)(220),
      output(25) => mem_array(25)(220),
      output(26) => mem_array(26)(220),
      output(27) => mem_array(27)(220),
      output(28) => mem_array(28)(220),
      output(29) => mem_array(29)(220),
      output(30) => mem_array(30)(220),
      output(31) => mem_array(31)(220),
      output(32) => mem_array(32)(220),
      output(33) => mem_array(33)(220),
      output(34) => mem_array(34)(220),
      output(35) => mem_array(35)(220)
      );
  rom221 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(221),
      output(0)  => mem_array(0)(221),
      output(1)  => mem_array(1)(221),
      output(2)  => mem_array(2)(221),
      output(3)  => mem_array(3)(221),
      output(4)  => mem_array(4)(221),
      output(5)  => mem_array(5)(221),
      output(6)  => mem_array(6)(221),
      output(7)  => mem_array(7)(221),
      output(8)  => mem_array(8)(221),
      output(9)  => mem_array(9)(221),
      output(10) => mem_array(10)(221),
      output(11) => mem_array(11)(221),
      output(12) => mem_array(12)(221),
      output(13) => mem_array(13)(221),
      output(14) => mem_array(14)(221),
      output(15) => mem_array(15)(221),
      output(16) => mem_array(16)(221),
      output(17) => mem_array(17)(221),
      output(18) => mem_array(18)(221),
      output(19) => mem_array(19)(221),
      output(20) => mem_array(20)(221),
      output(21) => mem_array(21)(221),
      output(22) => mem_array(22)(221),
      output(23) => mem_array(23)(221),
      output(24) => mem_array(24)(221),
      output(25) => mem_array(25)(221),
      output(26) => mem_array(26)(221),
      output(27) => mem_array(27)(221),
      output(28) => mem_array(28)(221),
      output(29) => mem_array(29)(221),
      output(30) => mem_array(30)(221),
      output(31) => mem_array(31)(221),
      output(32) => mem_array(32)(221),
      output(33) => mem_array(33)(221),
      output(34) => mem_array(34)(221),
      output(35) => mem_array(35)(221)
      );
  rom222 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(222),
      output(0)  => mem_array(0)(222),
      output(1)  => mem_array(1)(222),
      output(2)  => mem_array(2)(222),
      output(3)  => mem_array(3)(222),
      output(4)  => mem_array(4)(222),
      output(5)  => mem_array(5)(222),
      output(6)  => mem_array(6)(222),
      output(7)  => mem_array(7)(222),
      output(8)  => mem_array(8)(222),
      output(9)  => mem_array(9)(222),
      output(10) => mem_array(10)(222),
      output(11) => mem_array(11)(222),
      output(12) => mem_array(12)(222),
      output(13) => mem_array(13)(222),
      output(14) => mem_array(14)(222),
      output(15) => mem_array(15)(222),
      output(16) => mem_array(16)(222),
      output(17) => mem_array(17)(222),
      output(18) => mem_array(18)(222),
      output(19) => mem_array(19)(222),
      output(20) => mem_array(20)(222),
      output(21) => mem_array(21)(222),
      output(22) => mem_array(22)(222),
      output(23) => mem_array(23)(222),
      output(24) => mem_array(24)(222),
      output(25) => mem_array(25)(222),
      output(26) => mem_array(26)(222),
      output(27) => mem_array(27)(222),
      output(28) => mem_array(28)(222),
      output(29) => mem_array(29)(222),
      output(30) => mem_array(30)(222),
      output(31) => mem_array(31)(222),
      output(32) => mem_array(32)(222),
      output(33) => mem_array(33)(222),
      output(34) => mem_array(34)(222),
      output(35) => mem_array(35)(222)
      );
  rom223 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(223),
      output(0)  => mem_array(0)(223),
      output(1)  => mem_array(1)(223),
      output(2)  => mem_array(2)(223),
      output(3)  => mem_array(3)(223),
      output(4)  => mem_array(4)(223),
      output(5)  => mem_array(5)(223),
      output(6)  => mem_array(6)(223),
      output(7)  => mem_array(7)(223),
      output(8)  => mem_array(8)(223),
      output(9)  => mem_array(9)(223),
      output(10) => mem_array(10)(223),
      output(11) => mem_array(11)(223),
      output(12) => mem_array(12)(223),
      output(13) => mem_array(13)(223),
      output(14) => mem_array(14)(223),
      output(15) => mem_array(15)(223),
      output(16) => mem_array(16)(223),
      output(17) => mem_array(17)(223),
      output(18) => mem_array(18)(223),
      output(19) => mem_array(19)(223),
      output(20) => mem_array(20)(223),
      output(21) => mem_array(21)(223),
      output(22) => mem_array(22)(223),
      output(23) => mem_array(23)(223),
      output(24) => mem_array(24)(223),
      output(25) => mem_array(25)(223),
      output(26) => mem_array(26)(223),
      output(27) => mem_array(27)(223),
      output(28) => mem_array(28)(223),
      output(29) => mem_array(29)(223),
      output(30) => mem_array(30)(223),
      output(31) => mem_array(31)(223),
      output(32) => mem_array(32)(223),
      output(33) => mem_array(33)(223),
      output(34) => mem_array(34)(223),
      output(35) => mem_array(35)(223)
      );
  rom224 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(224),
      output(0)  => mem_array(0)(224),
      output(1)  => mem_array(1)(224),
      output(2)  => mem_array(2)(224),
      output(3)  => mem_array(3)(224),
      output(4)  => mem_array(4)(224),
      output(5)  => mem_array(5)(224),
      output(6)  => mem_array(6)(224),
      output(7)  => mem_array(7)(224),
      output(8)  => mem_array(8)(224),
      output(9)  => mem_array(9)(224),
      output(10) => mem_array(10)(224),
      output(11) => mem_array(11)(224),
      output(12) => mem_array(12)(224),
      output(13) => mem_array(13)(224),
      output(14) => mem_array(14)(224),
      output(15) => mem_array(15)(224),
      output(16) => mem_array(16)(224),
      output(17) => mem_array(17)(224),
      output(18) => mem_array(18)(224),
      output(19) => mem_array(19)(224),
      output(20) => mem_array(20)(224),
      output(21) => mem_array(21)(224),
      output(22) => mem_array(22)(224),
      output(23) => mem_array(23)(224),
      output(24) => mem_array(24)(224),
      output(25) => mem_array(25)(224),
      output(26) => mem_array(26)(224),
      output(27) => mem_array(27)(224),
      output(28) => mem_array(28)(224),
      output(29) => mem_array(29)(224),
      output(30) => mem_array(30)(224),
      output(31) => mem_array(31)(224),
      output(32) => mem_array(32)(224),
      output(33) => mem_array(33)(224),
      output(34) => mem_array(34)(224),
      output(35) => mem_array(35)(224)
      );
  rom225 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(225),
      output(0)  => mem_array(0)(225),
      output(1)  => mem_array(1)(225),
      output(2)  => mem_array(2)(225),
      output(3)  => mem_array(3)(225),
      output(4)  => mem_array(4)(225),
      output(5)  => mem_array(5)(225),
      output(6)  => mem_array(6)(225),
      output(7)  => mem_array(7)(225),
      output(8)  => mem_array(8)(225),
      output(9)  => mem_array(9)(225),
      output(10) => mem_array(10)(225),
      output(11) => mem_array(11)(225),
      output(12) => mem_array(12)(225),
      output(13) => mem_array(13)(225),
      output(14) => mem_array(14)(225),
      output(15) => mem_array(15)(225),
      output(16) => mem_array(16)(225),
      output(17) => mem_array(17)(225),
      output(18) => mem_array(18)(225),
      output(19) => mem_array(19)(225),
      output(20) => mem_array(20)(225),
      output(21) => mem_array(21)(225),
      output(22) => mem_array(22)(225),
      output(23) => mem_array(23)(225),
      output(24) => mem_array(24)(225),
      output(25) => mem_array(25)(225),
      output(26) => mem_array(26)(225),
      output(27) => mem_array(27)(225),
      output(28) => mem_array(28)(225),
      output(29) => mem_array(29)(225),
      output(30) => mem_array(30)(225),
      output(31) => mem_array(31)(225),
      output(32) => mem_array(32)(225),
      output(33) => mem_array(33)(225),
      output(34) => mem_array(34)(225),
      output(35) => mem_array(35)(225)
      );
  rom226 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(226),
      output(0)  => mem_array(0)(226),
      output(1)  => mem_array(1)(226),
      output(2)  => mem_array(2)(226),
      output(3)  => mem_array(3)(226),
      output(4)  => mem_array(4)(226),
      output(5)  => mem_array(5)(226),
      output(6)  => mem_array(6)(226),
      output(7)  => mem_array(7)(226),
      output(8)  => mem_array(8)(226),
      output(9)  => mem_array(9)(226),
      output(10) => mem_array(10)(226),
      output(11) => mem_array(11)(226),
      output(12) => mem_array(12)(226),
      output(13) => mem_array(13)(226),
      output(14) => mem_array(14)(226),
      output(15) => mem_array(15)(226),
      output(16) => mem_array(16)(226),
      output(17) => mem_array(17)(226),
      output(18) => mem_array(18)(226),
      output(19) => mem_array(19)(226),
      output(20) => mem_array(20)(226),
      output(21) => mem_array(21)(226),
      output(22) => mem_array(22)(226),
      output(23) => mem_array(23)(226),
      output(24) => mem_array(24)(226),
      output(25) => mem_array(25)(226),
      output(26) => mem_array(26)(226),
      output(27) => mem_array(27)(226),
      output(28) => mem_array(28)(226),
      output(29) => mem_array(29)(226),
      output(30) => mem_array(30)(226),
      output(31) => mem_array(31)(226),
      output(32) => mem_array(32)(226),
      output(33) => mem_array(33)(226),
      output(34) => mem_array(34)(226),
      output(35) => mem_array(35)(226)
      );
  rom227 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(227),
      output(0)  => mem_array(0)(227),
      output(1)  => mem_array(1)(227),
      output(2)  => mem_array(2)(227),
      output(3)  => mem_array(3)(227),
      output(4)  => mem_array(4)(227),
      output(5)  => mem_array(5)(227),
      output(6)  => mem_array(6)(227),
      output(7)  => mem_array(7)(227),
      output(8)  => mem_array(8)(227),
      output(9)  => mem_array(9)(227),
      output(10) => mem_array(10)(227),
      output(11) => mem_array(11)(227),
      output(12) => mem_array(12)(227),
      output(13) => mem_array(13)(227),
      output(14) => mem_array(14)(227),
      output(15) => mem_array(15)(227),
      output(16) => mem_array(16)(227),
      output(17) => mem_array(17)(227),
      output(18) => mem_array(18)(227),
      output(19) => mem_array(19)(227),
      output(20) => mem_array(20)(227),
      output(21) => mem_array(21)(227),
      output(22) => mem_array(22)(227),
      output(23) => mem_array(23)(227),
      output(24) => mem_array(24)(227),
      output(25) => mem_array(25)(227),
      output(26) => mem_array(26)(227),
      output(27) => mem_array(27)(227),
      output(28) => mem_array(28)(227),
      output(29) => mem_array(29)(227),
      output(30) => mem_array(30)(227),
      output(31) => mem_array(31)(227),
      output(32) => mem_array(32)(227),
      output(33) => mem_array(33)(227),
      output(34) => mem_array(34)(227),
      output(35) => mem_array(35)(227)
      );
  rom228 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(228),
      output(0)  => mem_array(0)(228),
      output(1)  => mem_array(1)(228),
      output(2)  => mem_array(2)(228),
      output(3)  => mem_array(3)(228),
      output(4)  => mem_array(4)(228),
      output(5)  => mem_array(5)(228),
      output(6)  => mem_array(6)(228),
      output(7)  => mem_array(7)(228),
      output(8)  => mem_array(8)(228),
      output(9)  => mem_array(9)(228),
      output(10) => mem_array(10)(228),
      output(11) => mem_array(11)(228),
      output(12) => mem_array(12)(228),
      output(13) => mem_array(13)(228),
      output(14) => mem_array(14)(228),
      output(15) => mem_array(15)(228),
      output(16) => mem_array(16)(228),
      output(17) => mem_array(17)(228),
      output(18) => mem_array(18)(228),
      output(19) => mem_array(19)(228),
      output(20) => mem_array(20)(228),
      output(21) => mem_array(21)(228),
      output(22) => mem_array(22)(228),
      output(23) => mem_array(23)(228),
      output(24) => mem_array(24)(228),
      output(25) => mem_array(25)(228),
      output(26) => mem_array(26)(228),
      output(27) => mem_array(27)(228),
      output(28) => mem_array(28)(228),
      output(29) => mem_array(29)(228),
      output(30) => mem_array(30)(228),
      output(31) => mem_array(31)(228),
      output(32) => mem_array(32)(228),
      output(33) => mem_array(33)(228),
      output(34) => mem_array(34)(228),
      output(35) => mem_array(35)(228)
      );
  rom229 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(229),
      output(0)  => mem_array(0)(229),
      output(1)  => mem_array(1)(229),
      output(2)  => mem_array(2)(229),
      output(3)  => mem_array(3)(229),
      output(4)  => mem_array(4)(229),
      output(5)  => mem_array(5)(229),
      output(6)  => mem_array(6)(229),
      output(7)  => mem_array(7)(229),
      output(8)  => mem_array(8)(229),
      output(9)  => mem_array(9)(229),
      output(10) => mem_array(10)(229),
      output(11) => mem_array(11)(229),
      output(12) => mem_array(12)(229),
      output(13) => mem_array(13)(229),
      output(14) => mem_array(14)(229),
      output(15) => mem_array(15)(229),
      output(16) => mem_array(16)(229),
      output(17) => mem_array(17)(229),
      output(18) => mem_array(18)(229),
      output(19) => mem_array(19)(229),
      output(20) => mem_array(20)(229),
      output(21) => mem_array(21)(229),
      output(22) => mem_array(22)(229),
      output(23) => mem_array(23)(229),
      output(24) => mem_array(24)(229),
      output(25) => mem_array(25)(229),
      output(26) => mem_array(26)(229),
      output(27) => mem_array(27)(229),
      output(28) => mem_array(28)(229),
      output(29) => mem_array(29)(229),
      output(30) => mem_array(30)(229),
      output(31) => mem_array(31)(229),
      output(32) => mem_array(32)(229),
      output(33) => mem_array(33)(229),
      output(34) => mem_array(34)(229),
      output(35) => mem_array(35)(229)
      );
  rom230 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(230),
      output(0)  => mem_array(0)(230),
      output(1)  => mem_array(1)(230),
      output(2)  => mem_array(2)(230),
      output(3)  => mem_array(3)(230),
      output(4)  => mem_array(4)(230),
      output(5)  => mem_array(5)(230),
      output(6)  => mem_array(6)(230),
      output(7)  => mem_array(7)(230),
      output(8)  => mem_array(8)(230),
      output(9)  => mem_array(9)(230),
      output(10) => mem_array(10)(230),
      output(11) => mem_array(11)(230),
      output(12) => mem_array(12)(230),
      output(13) => mem_array(13)(230),
      output(14) => mem_array(14)(230),
      output(15) => mem_array(15)(230),
      output(16) => mem_array(16)(230),
      output(17) => mem_array(17)(230),
      output(18) => mem_array(18)(230),
      output(19) => mem_array(19)(230),
      output(20) => mem_array(20)(230),
      output(21) => mem_array(21)(230),
      output(22) => mem_array(22)(230),
      output(23) => mem_array(23)(230),
      output(24) => mem_array(24)(230),
      output(25) => mem_array(25)(230),
      output(26) => mem_array(26)(230),
      output(27) => mem_array(27)(230),
      output(28) => mem_array(28)(230),
      output(29) => mem_array(29)(230),
      output(30) => mem_array(30)(230),
      output(31) => mem_array(31)(230),
      output(32) => mem_array(32)(230),
      output(33) => mem_array(33)(230),
      output(34) => mem_array(34)(230),
      output(35) => mem_array(35)(230)
      );
  rom231 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(231),
      output(0)  => mem_array(0)(231),
      output(1)  => mem_array(1)(231),
      output(2)  => mem_array(2)(231),
      output(3)  => mem_array(3)(231),
      output(4)  => mem_array(4)(231),
      output(5)  => mem_array(5)(231),
      output(6)  => mem_array(6)(231),
      output(7)  => mem_array(7)(231),
      output(8)  => mem_array(8)(231),
      output(9)  => mem_array(9)(231),
      output(10) => mem_array(10)(231),
      output(11) => mem_array(11)(231),
      output(12) => mem_array(12)(231),
      output(13) => mem_array(13)(231),
      output(14) => mem_array(14)(231),
      output(15) => mem_array(15)(231),
      output(16) => mem_array(16)(231),
      output(17) => mem_array(17)(231),
      output(18) => mem_array(18)(231),
      output(19) => mem_array(19)(231),
      output(20) => mem_array(20)(231),
      output(21) => mem_array(21)(231),
      output(22) => mem_array(22)(231),
      output(23) => mem_array(23)(231),
      output(24) => mem_array(24)(231),
      output(25) => mem_array(25)(231),
      output(26) => mem_array(26)(231),
      output(27) => mem_array(27)(231),
      output(28) => mem_array(28)(231),
      output(29) => mem_array(29)(231),
      output(30) => mem_array(30)(231),
      output(31) => mem_array(31)(231),
      output(32) => mem_array(32)(231),
      output(33) => mem_array(33)(231),
      output(34) => mem_array(34)(231),
      output(35) => mem_array(35)(231)
      );
  rom232 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(232),
      output(0)  => mem_array(0)(232),
      output(1)  => mem_array(1)(232),
      output(2)  => mem_array(2)(232),
      output(3)  => mem_array(3)(232),
      output(4)  => mem_array(4)(232),
      output(5)  => mem_array(5)(232),
      output(6)  => mem_array(6)(232),
      output(7)  => mem_array(7)(232),
      output(8)  => mem_array(8)(232),
      output(9)  => mem_array(9)(232),
      output(10) => mem_array(10)(232),
      output(11) => mem_array(11)(232),
      output(12) => mem_array(12)(232),
      output(13) => mem_array(13)(232),
      output(14) => mem_array(14)(232),
      output(15) => mem_array(15)(232),
      output(16) => mem_array(16)(232),
      output(17) => mem_array(17)(232),
      output(18) => mem_array(18)(232),
      output(19) => mem_array(19)(232),
      output(20) => mem_array(20)(232),
      output(21) => mem_array(21)(232),
      output(22) => mem_array(22)(232),
      output(23) => mem_array(23)(232),
      output(24) => mem_array(24)(232),
      output(25) => mem_array(25)(232),
      output(26) => mem_array(26)(232),
      output(27) => mem_array(27)(232),
      output(28) => mem_array(28)(232),
      output(29) => mem_array(29)(232),
      output(30) => mem_array(30)(232),
      output(31) => mem_array(31)(232),
      output(32) => mem_array(32)(232),
      output(33) => mem_array(33)(232),
      output(34) => mem_array(34)(232),
      output(35) => mem_array(35)(232)
      );
  rom233 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(233),
      output(0)  => mem_array(0)(233),
      output(1)  => mem_array(1)(233),
      output(2)  => mem_array(2)(233),
      output(3)  => mem_array(3)(233),
      output(4)  => mem_array(4)(233),
      output(5)  => mem_array(5)(233),
      output(6)  => mem_array(6)(233),
      output(7)  => mem_array(7)(233),
      output(8)  => mem_array(8)(233),
      output(9)  => mem_array(9)(233),
      output(10) => mem_array(10)(233),
      output(11) => mem_array(11)(233),
      output(12) => mem_array(12)(233),
      output(13) => mem_array(13)(233),
      output(14) => mem_array(14)(233),
      output(15) => mem_array(15)(233),
      output(16) => mem_array(16)(233),
      output(17) => mem_array(17)(233),
      output(18) => mem_array(18)(233),
      output(19) => mem_array(19)(233),
      output(20) => mem_array(20)(233),
      output(21) => mem_array(21)(233),
      output(22) => mem_array(22)(233),
      output(23) => mem_array(23)(233),
      output(24) => mem_array(24)(233),
      output(25) => mem_array(25)(233),
      output(26) => mem_array(26)(233),
      output(27) => mem_array(27)(233),
      output(28) => mem_array(28)(233),
      output(29) => mem_array(29)(233),
      output(30) => mem_array(30)(233),
      output(31) => mem_array(31)(233),
      output(32) => mem_array(32)(233),
      output(33) => mem_array(33)(233),
      output(34) => mem_array(34)(233),
      output(35) => mem_array(35)(233)
      );
  rom234 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(234),
      output(0)  => mem_array(0)(234),
      output(1)  => mem_array(1)(234),
      output(2)  => mem_array(2)(234),
      output(3)  => mem_array(3)(234),
      output(4)  => mem_array(4)(234),
      output(5)  => mem_array(5)(234),
      output(6)  => mem_array(6)(234),
      output(7)  => mem_array(7)(234),
      output(8)  => mem_array(8)(234),
      output(9)  => mem_array(9)(234),
      output(10) => mem_array(10)(234),
      output(11) => mem_array(11)(234),
      output(12) => mem_array(12)(234),
      output(13) => mem_array(13)(234),
      output(14) => mem_array(14)(234),
      output(15) => mem_array(15)(234),
      output(16) => mem_array(16)(234),
      output(17) => mem_array(17)(234),
      output(18) => mem_array(18)(234),
      output(19) => mem_array(19)(234),
      output(20) => mem_array(20)(234),
      output(21) => mem_array(21)(234),
      output(22) => mem_array(22)(234),
      output(23) => mem_array(23)(234),
      output(24) => mem_array(24)(234),
      output(25) => mem_array(25)(234),
      output(26) => mem_array(26)(234),
      output(27) => mem_array(27)(234),
      output(28) => mem_array(28)(234),
      output(29) => mem_array(29)(234),
      output(30) => mem_array(30)(234),
      output(31) => mem_array(31)(234),
      output(32) => mem_array(32)(234),
      output(33) => mem_array(33)(234),
      output(34) => mem_array(34)(234),
      output(35) => mem_array(35)(234)
      );
  rom235 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(235),
      output(0)  => mem_array(0)(235),
      output(1)  => mem_array(1)(235),
      output(2)  => mem_array(2)(235),
      output(3)  => mem_array(3)(235),
      output(4)  => mem_array(4)(235),
      output(5)  => mem_array(5)(235),
      output(6)  => mem_array(6)(235),
      output(7)  => mem_array(7)(235),
      output(8)  => mem_array(8)(235),
      output(9)  => mem_array(9)(235),
      output(10) => mem_array(10)(235),
      output(11) => mem_array(11)(235),
      output(12) => mem_array(12)(235),
      output(13) => mem_array(13)(235),
      output(14) => mem_array(14)(235),
      output(15) => mem_array(15)(235),
      output(16) => mem_array(16)(235),
      output(17) => mem_array(17)(235),
      output(18) => mem_array(18)(235),
      output(19) => mem_array(19)(235),
      output(20) => mem_array(20)(235),
      output(21) => mem_array(21)(235),
      output(22) => mem_array(22)(235),
      output(23) => mem_array(23)(235),
      output(24) => mem_array(24)(235),
      output(25) => mem_array(25)(235),
      output(26) => mem_array(26)(235),
      output(27) => mem_array(27)(235),
      output(28) => mem_array(28)(235),
      output(29) => mem_array(29)(235),
      output(30) => mem_array(30)(235),
      output(31) => mem_array(31)(235),
      output(32) => mem_array(32)(235),
      output(33) => mem_array(33)(235),
      output(34) => mem_array(34)(235),
      output(35) => mem_array(35)(235)
      );
  rom236 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(236),
      output(0)  => mem_array(0)(236),
      output(1)  => mem_array(1)(236),
      output(2)  => mem_array(2)(236),
      output(3)  => mem_array(3)(236),
      output(4)  => mem_array(4)(236),
      output(5)  => mem_array(5)(236),
      output(6)  => mem_array(6)(236),
      output(7)  => mem_array(7)(236),
      output(8)  => mem_array(8)(236),
      output(9)  => mem_array(9)(236),
      output(10) => mem_array(10)(236),
      output(11) => mem_array(11)(236),
      output(12) => mem_array(12)(236),
      output(13) => mem_array(13)(236),
      output(14) => mem_array(14)(236),
      output(15) => mem_array(15)(236),
      output(16) => mem_array(16)(236),
      output(17) => mem_array(17)(236),
      output(18) => mem_array(18)(236),
      output(19) => mem_array(19)(236),
      output(20) => mem_array(20)(236),
      output(21) => mem_array(21)(236),
      output(22) => mem_array(22)(236),
      output(23) => mem_array(23)(236),
      output(24) => mem_array(24)(236),
      output(25) => mem_array(25)(236),
      output(26) => mem_array(26)(236),
      output(27) => mem_array(27)(236),
      output(28) => mem_array(28)(236),
      output(29) => mem_array(29)(236),
      output(30) => mem_array(30)(236),
      output(31) => mem_array(31)(236),
      output(32) => mem_array(32)(236),
      output(33) => mem_array(33)(236),
      output(34) => mem_array(34)(236),
      output(35) => mem_array(35)(236)
      );
  rom237 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(237),
      output(0)  => mem_array(0)(237),
      output(1)  => mem_array(1)(237),
      output(2)  => mem_array(2)(237),
      output(3)  => mem_array(3)(237),
      output(4)  => mem_array(4)(237),
      output(5)  => mem_array(5)(237),
      output(6)  => mem_array(6)(237),
      output(7)  => mem_array(7)(237),
      output(8)  => mem_array(8)(237),
      output(9)  => mem_array(9)(237),
      output(10) => mem_array(10)(237),
      output(11) => mem_array(11)(237),
      output(12) => mem_array(12)(237),
      output(13) => mem_array(13)(237),
      output(14) => mem_array(14)(237),
      output(15) => mem_array(15)(237),
      output(16) => mem_array(16)(237),
      output(17) => mem_array(17)(237),
      output(18) => mem_array(18)(237),
      output(19) => mem_array(19)(237),
      output(20) => mem_array(20)(237),
      output(21) => mem_array(21)(237),
      output(22) => mem_array(22)(237),
      output(23) => mem_array(23)(237),
      output(24) => mem_array(24)(237),
      output(25) => mem_array(25)(237),
      output(26) => mem_array(26)(237),
      output(27) => mem_array(27)(237),
      output(28) => mem_array(28)(237),
      output(29) => mem_array(29)(237),
      output(30) => mem_array(30)(237),
      output(31) => mem_array(31)(237),
      output(32) => mem_array(32)(237),
      output(33) => mem_array(33)(237),
      output(34) => mem_array(34)(237),
      output(35) => mem_array(35)(237)
      );
  rom238 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(238),
      output(0)  => mem_array(0)(238),
      output(1)  => mem_array(1)(238),
      output(2)  => mem_array(2)(238),
      output(3)  => mem_array(3)(238),
      output(4)  => mem_array(4)(238),
      output(5)  => mem_array(5)(238),
      output(6)  => mem_array(6)(238),
      output(7)  => mem_array(7)(238),
      output(8)  => mem_array(8)(238),
      output(9)  => mem_array(9)(238),
      output(10) => mem_array(10)(238),
      output(11) => mem_array(11)(238),
      output(12) => mem_array(12)(238),
      output(13) => mem_array(13)(238),
      output(14) => mem_array(14)(238),
      output(15) => mem_array(15)(238),
      output(16) => mem_array(16)(238),
      output(17) => mem_array(17)(238),
      output(18) => mem_array(18)(238),
      output(19) => mem_array(19)(238),
      output(20) => mem_array(20)(238),
      output(21) => mem_array(21)(238),
      output(22) => mem_array(22)(238),
      output(23) => mem_array(23)(238),
      output(24) => mem_array(24)(238),
      output(25) => mem_array(25)(238),
      output(26) => mem_array(26)(238),
      output(27) => mem_array(27)(238),
      output(28) => mem_array(28)(238),
      output(29) => mem_array(29)(238),
      output(30) => mem_array(30)(238),
      output(31) => mem_array(31)(238),
      output(32) => mem_array(32)(238),
      output(33) => mem_array(33)(238),
      output(34) => mem_array(34)(238),
      output(35) => mem_array(35)(238)
      );
  rom239 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(239),
      output(0)  => mem_array(0)(239),
      output(1)  => mem_array(1)(239),
      output(2)  => mem_array(2)(239),
      output(3)  => mem_array(3)(239),
      output(4)  => mem_array(4)(239),
      output(5)  => mem_array(5)(239),
      output(6)  => mem_array(6)(239),
      output(7)  => mem_array(7)(239),
      output(8)  => mem_array(8)(239),
      output(9)  => mem_array(9)(239),
      output(10) => mem_array(10)(239),
      output(11) => mem_array(11)(239),
      output(12) => mem_array(12)(239),
      output(13) => mem_array(13)(239),
      output(14) => mem_array(14)(239),
      output(15) => mem_array(15)(239),
      output(16) => mem_array(16)(239),
      output(17) => mem_array(17)(239),
      output(18) => mem_array(18)(239),
      output(19) => mem_array(19)(239),
      output(20) => mem_array(20)(239),
      output(21) => mem_array(21)(239),
      output(22) => mem_array(22)(239),
      output(23) => mem_array(23)(239),
      output(24) => mem_array(24)(239),
      output(25) => mem_array(25)(239),
      output(26) => mem_array(26)(239),
      output(27) => mem_array(27)(239),
      output(28) => mem_array(28)(239),
      output(29) => mem_array(29)(239),
      output(30) => mem_array(30)(239),
      output(31) => mem_array(31)(239),
      output(32) => mem_array(32)(239),
      output(33) => mem_array(33)(239),
      output(34) => mem_array(34)(239),
      output(35) => mem_array(35)(239)
      );
  rom240 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(240),
      output(0)  => mem_array(0)(240),
      output(1)  => mem_array(1)(240),
      output(2)  => mem_array(2)(240),
      output(3)  => mem_array(3)(240),
      output(4)  => mem_array(4)(240),
      output(5)  => mem_array(5)(240),
      output(6)  => mem_array(6)(240),
      output(7)  => mem_array(7)(240),
      output(8)  => mem_array(8)(240),
      output(9)  => mem_array(9)(240),
      output(10) => mem_array(10)(240),
      output(11) => mem_array(11)(240),
      output(12) => mem_array(12)(240),
      output(13) => mem_array(13)(240),
      output(14) => mem_array(14)(240),
      output(15) => mem_array(15)(240),
      output(16) => mem_array(16)(240),
      output(17) => mem_array(17)(240),
      output(18) => mem_array(18)(240),
      output(19) => mem_array(19)(240),
      output(20) => mem_array(20)(240),
      output(21) => mem_array(21)(240),
      output(22) => mem_array(22)(240),
      output(23) => mem_array(23)(240),
      output(24) => mem_array(24)(240),
      output(25) => mem_array(25)(240),
      output(26) => mem_array(26)(240),
      output(27) => mem_array(27)(240),
      output(28) => mem_array(28)(240),
      output(29) => mem_array(29)(240),
      output(30) => mem_array(30)(240),
      output(31) => mem_array(31)(240),
      output(32) => mem_array(32)(240),
      output(33) => mem_array(33)(240),
      output(34) => mem_array(34)(240),
      output(35) => mem_array(35)(240)
      );
  rom241 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(241),
      output(0)  => mem_array(0)(241),
      output(1)  => mem_array(1)(241),
      output(2)  => mem_array(2)(241),
      output(3)  => mem_array(3)(241),
      output(4)  => mem_array(4)(241),
      output(5)  => mem_array(5)(241),
      output(6)  => mem_array(6)(241),
      output(7)  => mem_array(7)(241),
      output(8)  => mem_array(8)(241),
      output(9)  => mem_array(9)(241),
      output(10) => mem_array(10)(241),
      output(11) => mem_array(11)(241),
      output(12) => mem_array(12)(241),
      output(13) => mem_array(13)(241),
      output(14) => mem_array(14)(241),
      output(15) => mem_array(15)(241),
      output(16) => mem_array(16)(241),
      output(17) => mem_array(17)(241),
      output(18) => mem_array(18)(241),
      output(19) => mem_array(19)(241),
      output(20) => mem_array(20)(241),
      output(21) => mem_array(21)(241),
      output(22) => mem_array(22)(241),
      output(23) => mem_array(23)(241),
      output(24) => mem_array(24)(241),
      output(25) => mem_array(25)(241),
      output(26) => mem_array(26)(241),
      output(27) => mem_array(27)(241),
      output(28) => mem_array(28)(241),
      output(29) => mem_array(29)(241),
      output(30) => mem_array(30)(241),
      output(31) => mem_array(31)(241),
      output(32) => mem_array(32)(241),
      output(33) => mem_array(33)(241),
      output(34) => mem_array(34)(241),
      output(35) => mem_array(35)(241)
      );
  rom242 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(242),
      output(0)  => mem_array(0)(242),
      output(1)  => mem_array(1)(242),
      output(2)  => mem_array(2)(242),
      output(3)  => mem_array(3)(242),
      output(4)  => mem_array(4)(242),
      output(5)  => mem_array(5)(242),
      output(6)  => mem_array(6)(242),
      output(7)  => mem_array(7)(242),
      output(8)  => mem_array(8)(242),
      output(9)  => mem_array(9)(242),
      output(10) => mem_array(10)(242),
      output(11) => mem_array(11)(242),
      output(12) => mem_array(12)(242),
      output(13) => mem_array(13)(242),
      output(14) => mem_array(14)(242),
      output(15) => mem_array(15)(242),
      output(16) => mem_array(16)(242),
      output(17) => mem_array(17)(242),
      output(18) => mem_array(18)(242),
      output(19) => mem_array(19)(242),
      output(20) => mem_array(20)(242),
      output(21) => mem_array(21)(242),
      output(22) => mem_array(22)(242),
      output(23) => mem_array(23)(242),
      output(24) => mem_array(24)(242),
      output(25) => mem_array(25)(242),
      output(26) => mem_array(26)(242),
      output(27) => mem_array(27)(242),
      output(28) => mem_array(28)(242),
      output(29) => mem_array(29)(242),
      output(30) => mem_array(30)(242),
      output(31) => mem_array(31)(242),
      output(32) => mem_array(32)(242),
      output(33) => mem_array(33)(242),
      output(34) => mem_array(34)(242),
      output(35) => mem_array(35)(242)
      );
  rom243 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(243),
      output(0)  => mem_array(0)(243),
      output(1)  => mem_array(1)(243),
      output(2)  => mem_array(2)(243),
      output(3)  => mem_array(3)(243),
      output(4)  => mem_array(4)(243),
      output(5)  => mem_array(5)(243),
      output(6)  => mem_array(6)(243),
      output(7)  => mem_array(7)(243),
      output(8)  => mem_array(8)(243),
      output(9)  => mem_array(9)(243),
      output(10) => mem_array(10)(243),
      output(11) => mem_array(11)(243),
      output(12) => mem_array(12)(243),
      output(13) => mem_array(13)(243),
      output(14) => mem_array(14)(243),
      output(15) => mem_array(15)(243),
      output(16) => mem_array(16)(243),
      output(17) => mem_array(17)(243),
      output(18) => mem_array(18)(243),
      output(19) => mem_array(19)(243),
      output(20) => mem_array(20)(243),
      output(21) => mem_array(21)(243),
      output(22) => mem_array(22)(243),
      output(23) => mem_array(23)(243),
      output(24) => mem_array(24)(243),
      output(25) => mem_array(25)(243),
      output(26) => mem_array(26)(243),
      output(27) => mem_array(27)(243),
      output(28) => mem_array(28)(243),
      output(29) => mem_array(29)(243),
      output(30) => mem_array(30)(243),
      output(31) => mem_array(31)(243),
      output(32) => mem_array(32)(243),
      output(33) => mem_array(33)(243),
      output(34) => mem_array(34)(243),
      output(35) => mem_array(35)(243)
      );
  rom244 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(244),
      output(0)  => mem_array(0)(244),
      output(1)  => mem_array(1)(244),
      output(2)  => mem_array(2)(244),
      output(3)  => mem_array(3)(244),
      output(4)  => mem_array(4)(244),
      output(5)  => mem_array(5)(244),
      output(6)  => mem_array(6)(244),
      output(7)  => mem_array(7)(244),
      output(8)  => mem_array(8)(244),
      output(9)  => mem_array(9)(244),
      output(10) => mem_array(10)(244),
      output(11) => mem_array(11)(244),
      output(12) => mem_array(12)(244),
      output(13) => mem_array(13)(244),
      output(14) => mem_array(14)(244),
      output(15) => mem_array(15)(244),
      output(16) => mem_array(16)(244),
      output(17) => mem_array(17)(244),
      output(18) => mem_array(18)(244),
      output(19) => mem_array(19)(244),
      output(20) => mem_array(20)(244),
      output(21) => mem_array(21)(244),
      output(22) => mem_array(22)(244),
      output(23) => mem_array(23)(244),
      output(24) => mem_array(24)(244),
      output(25) => mem_array(25)(244),
      output(26) => mem_array(26)(244),
      output(27) => mem_array(27)(244),
      output(28) => mem_array(28)(244),
      output(29) => mem_array(29)(244),
      output(30) => mem_array(30)(244),
      output(31) => mem_array(31)(244),
      output(32) => mem_array(32)(244),
      output(33) => mem_array(33)(244),
      output(34) => mem_array(34)(244),
      output(35) => mem_array(35)(244)
      );
  rom245 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(245),
      output(0)  => mem_array(0)(245),
      output(1)  => mem_array(1)(245),
      output(2)  => mem_array(2)(245),
      output(3)  => mem_array(3)(245),
      output(4)  => mem_array(4)(245),
      output(5)  => mem_array(5)(245),
      output(6)  => mem_array(6)(245),
      output(7)  => mem_array(7)(245),
      output(8)  => mem_array(8)(245),
      output(9)  => mem_array(9)(245),
      output(10) => mem_array(10)(245),
      output(11) => mem_array(11)(245),
      output(12) => mem_array(12)(245),
      output(13) => mem_array(13)(245),
      output(14) => mem_array(14)(245),
      output(15) => mem_array(15)(245),
      output(16) => mem_array(16)(245),
      output(17) => mem_array(17)(245),
      output(18) => mem_array(18)(245),
      output(19) => mem_array(19)(245),
      output(20) => mem_array(20)(245),
      output(21) => mem_array(21)(245),
      output(22) => mem_array(22)(245),
      output(23) => mem_array(23)(245),
      output(24) => mem_array(24)(245),
      output(25) => mem_array(25)(245),
      output(26) => mem_array(26)(245),
      output(27) => mem_array(27)(245),
      output(28) => mem_array(28)(245),
      output(29) => mem_array(29)(245),
      output(30) => mem_array(30)(245),
      output(31) => mem_array(31)(245),
      output(32) => mem_array(32)(245),
      output(33) => mem_array(33)(245),
      output(34) => mem_array(34)(245),
      output(35) => mem_array(35)(245)
      );
  rom246 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(246),
      output(0)  => mem_array(0)(246),
      output(1)  => mem_array(1)(246),
      output(2)  => mem_array(2)(246),
      output(3)  => mem_array(3)(246),
      output(4)  => mem_array(4)(246),
      output(5)  => mem_array(5)(246),
      output(6)  => mem_array(6)(246),
      output(7)  => mem_array(7)(246),
      output(8)  => mem_array(8)(246),
      output(9)  => mem_array(9)(246),
      output(10) => mem_array(10)(246),
      output(11) => mem_array(11)(246),
      output(12) => mem_array(12)(246),
      output(13) => mem_array(13)(246),
      output(14) => mem_array(14)(246),
      output(15) => mem_array(15)(246),
      output(16) => mem_array(16)(246),
      output(17) => mem_array(17)(246),
      output(18) => mem_array(18)(246),
      output(19) => mem_array(19)(246),
      output(20) => mem_array(20)(246),
      output(21) => mem_array(21)(246),
      output(22) => mem_array(22)(246),
      output(23) => mem_array(23)(246),
      output(24) => mem_array(24)(246),
      output(25) => mem_array(25)(246),
      output(26) => mem_array(26)(246),
      output(27) => mem_array(27)(246),
      output(28) => mem_array(28)(246),
      output(29) => mem_array(29)(246),
      output(30) => mem_array(30)(246),
      output(31) => mem_array(31)(246),
      output(32) => mem_array(32)(246),
      output(33) => mem_array(33)(246),
      output(34) => mem_array(34)(246),
      output(35) => mem_array(35)(246)
      );
  rom247 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(247),
      output(0)  => mem_array(0)(247),
      output(1)  => mem_array(1)(247),
      output(2)  => mem_array(2)(247),
      output(3)  => mem_array(3)(247),
      output(4)  => mem_array(4)(247),
      output(5)  => mem_array(5)(247),
      output(6)  => mem_array(6)(247),
      output(7)  => mem_array(7)(247),
      output(8)  => mem_array(8)(247),
      output(9)  => mem_array(9)(247),
      output(10) => mem_array(10)(247),
      output(11) => mem_array(11)(247),
      output(12) => mem_array(12)(247),
      output(13) => mem_array(13)(247),
      output(14) => mem_array(14)(247),
      output(15) => mem_array(15)(247),
      output(16) => mem_array(16)(247),
      output(17) => mem_array(17)(247),
      output(18) => mem_array(18)(247),
      output(19) => mem_array(19)(247),
      output(20) => mem_array(20)(247),
      output(21) => mem_array(21)(247),
      output(22) => mem_array(22)(247),
      output(23) => mem_array(23)(247),
      output(24) => mem_array(24)(247),
      output(25) => mem_array(25)(247),
      output(26) => mem_array(26)(247),
      output(27) => mem_array(27)(247),
      output(28) => mem_array(28)(247),
      output(29) => mem_array(29)(247),
      output(30) => mem_array(30)(247),
      output(31) => mem_array(31)(247),
      output(32) => mem_array(32)(247),
      output(33) => mem_array(33)(247),
      output(34) => mem_array(34)(247),
      output(35) => mem_array(35)(247)
      );
  rom248 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(248),
      output(0)  => mem_array(0)(248),
      output(1)  => mem_array(1)(248),
      output(2)  => mem_array(2)(248),
      output(3)  => mem_array(3)(248),
      output(4)  => mem_array(4)(248),
      output(5)  => mem_array(5)(248),
      output(6)  => mem_array(6)(248),
      output(7)  => mem_array(7)(248),
      output(8)  => mem_array(8)(248),
      output(9)  => mem_array(9)(248),
      output(10) => mem_array(10)(248),
      output(11) => mem_array(11)(248),
      output(12) => mem_array(12)(248),
      output(13) => mem_array(13)(248),
      output(14) => mem_array(14)(248),
      output(15) => mem_array(15)(248),
      output(16) => mem_array(16)(248),
      output(17) => mem_array(17)(248),
      output(18) => mem_array(18)(248),
      output(19) => mem_array(19)(248),
      output(20) => mem_array(20)(248),
      output(21) => mem_array(21)(248),
      output(22) => mem_array(22)(248),
      output(23) => mem_array(23)(248),
      output(24) => mem_array(24)(248),
      output(25) => mem_array(25)(248),
      output(26) => mem_array(26)(248),
      output(27) => mem_array(27)(248),
      output(28) => mem_array(28)(248),
      output(29) => mem_array(29)(248),
      output(30) => mem_array(30)(248),
      output(31) => mem_array(31)(248),
      output(32) => mem_array(32)(248),
      output(33) => mem_array(33)(248),
      output(34) => mem_array(34)(248),
      output(35) => mem_array(35)(248)
      );
  rom249 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(249),
      output(0)  => mem_array(0)(249),
      output(1)  => mem_array(1)(249),
      output(2)  => mem_array(2)(249),
      output(3)  => mem_array(3)(249),
      output(4)  => mem_array(4)(249),
      output(5)  => mem_array(5)(249),
      output(6)  => mem_array(6)(249),
      output(7)  => mem_array(7)(249),
      output(8)  => mem_array(8)(249),
      output(9)  => mem_array(9)(249),
      output(10) => mem_array(10)(249),
      output(11) => mem_array(11)(249),
      output(12) => mem_array(12)(249),
      output(13) => mem_array(13)(249),
      output(14) => mem_array(14)(249),
      output(15) => mem_array(15)(249),
      output(16) => mem_array(16)(249),
      output(17) => mem_array(17)(249),
      output(18) => mem_array(18)(249),
      output(19) => mem_array(19)(249),
      output(20) => mem_array(20)(249),
      output(21) => mem_array(21)(249),
      output(22) => mem_array(22)(249),
      output(23) => mem_array(23)(249),
      output(24) => mem_array(24)(249),
      output(25) => mem_array(25)(249),
      output(26) => mem_array(26)(249),
      output(27) => mem_array(27)(249),
      output(28) => mem_array(28)(249),
      output(29) => mem_array(29)(249),
      output(30) => mem_array(30)(249),
      output(31) => mem_array(31)(249),
      output(32) => mem_array(32)(249),
      output(33) => mem_array(33)(249),
      output(34) => mem_array(34)(249),
      output(35) => mem_array(35)(249)
      );
  rom250 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(250),
      output(0)  => mem_array(0)(250),
      output(1)  => mem_array(1)(250),
      output(2)  => mem_array(2)(250),
      output(3)  => mem_array(3)(250),
      output(4)  => mem_array(4)(250),
      output(5)  => mem_array(5)(250),
      output(6)  => mem_array(6)(250),
      output(7)  => mem_array(7)(250),
      output(8)  => mem_array(8)(250),
      output(9)  => mem_array(9)(250),
      output(10) => mem_array(10)(250),
      output(11) => mem_array(11)(250),
      output(12) => mem_array(12)(250),
      output(13) => mem_array(13)(250),
      output(14) => mem_array(14)(250),
      output(15) => mem_array(15)(250),
      output(16) => mem_array(16)(250),
      output(17) => mem_array(17)(250),
      output(18) => mem_array(18)(250),
      output(19) => mem_array(19)(250),
      output(20) => mem_array(20)(250),
      output(21) => mem_array(21)(250),
      output(22) => mem_array(22)(250),
      output(23) => mem_array(23)(250),
      output(24) => mem_array(24)(250),
      output(25) => mem_array(25)(250),
      output(26) => mem_array(26)(250),
      output(27) => mem_array(27)(250),
      output(28) => mem_array(28)(250),
      output(29) => mem_array(29)(250),
      output(30) => mem_array(30)(250),
      output(31) => mem_array(31)(250),
      output(32) => mem_array(32)(250),
      output(33) => mem_array(33)(250),
      output(34) => mem_array(34)(250),
      output(35) => mem_array(35)(250)
      );
  rom251 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(251),
      output(0)  => mem_array(0)(251),
      output(1)  => mem_array(1)(251),
      output(2)  => mem_array(2)(251),
      output(3)  => mem_array(3)(251),
      output(4)  => mem_array(4)(251),
      output(5)  => mem_array(5)(251),
      output(6)  => mem_array(6)(251),
      output(7)  => mem_array(7)(251),
      output(8)  => mem_array(8)(251),
      output(9)  => mem_array(9)(251),
      output(10) => mem_array(10)(251),
      output(11) => mem_array(11)(251),
      output(12) => mem_array(12)(251),
      output(13) => mem_array(13)(251),
      output(14) => mem_array(14)(251),
      output(15) => mem_array(15)(251),
      output(16) => mem_array(16)(251),
      output(17) => mem_array(17)(251),
      output(18) => mem_array(18)(251),
      output(19) => mem_array(19)(251),
      output(20) => mem_array(20)(251),
      output(21) => mem_array(21)(251),
      output(22) => mem_array(22)(251),
      output(23) => mem_array(23)(251),
      output(24) => mem_array(24)(251),
      output(25) => mem_array(25)(251),
      output(26) => mem_array(26)(251),
      output(27) => mem_array(27)(251),
      output(28) => mem_array(28)(251),
      output(29) => mem_array(29)(251),
      output(30) => mem_array(30)(251),
      output(31) => mem_array(31)(251),
      output(32) => mem_array(32)(251),
      output(33) => mem_array(33)(251),
      output(34) => mem_array(34)(251),
      output(35) => mem_array(35)(251)
      );
  rom252 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(252),
      output(0)  => mem_array(0)(252),
      output(1)  => mem_array(1)(252),
      output(2)  => mem_array(2)(252),
      output(3)  => mem_array(3)(252),
      output(4)  => mem_array(4)(252),
      output(5)  => mem_array(5)(252),
      output(6)  => mem_array(6)(252),
      output(7)  => mem_array(7)(252),
      output(8)  => mem_array(8)(252),
      output(9)  => mem_array(9)(252),
      output(10) => mem_array(10)(252),
      output(11) => mem_array(11)(252),
      output(12) => mem_array(12)(252),
      output(13) => mem_array(13)(252),
      output(14) => mem_array(14)(252),
      output(15) => mem_array(15)(252),
      output(16) => mem_array(16)(252),
      output(17) => mem_array(17)(252),
      output(18) => mem_array(18)(252),
      output(19) => mem_array(19)(252),
      output(20) => mem_array(20)(252),
      output(21) => mem_array(21)(252),
      output(22) => mem_array(22)(252),
      output(23) => mem_array(23)(252),
      output(24) => mem_array(24)(252),
      output(25) => mem_array(25)(252),
      output(26) => mem_array(26)(252),
      output(27) => mem_array(27)(252),
      output(28) => mem_array(28)(252),
      output(29) => mem_array(29)(252),
      output(30) => mem_array(30)(252),
      output(31) => mem_array(31)(252),
      output(32) => mem_array(32)(252),
      output(33) => mem_array(33)(252),
      output(34) => mem_array(34)(252),
      output(35) => mem_array(35)(252)
      );
  rom253 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(253),
      output(0)  => mem_array(0)(253),
      output(1)  => mem_array(1)(253),
      output(2)  => mem_array(2)(253),
      output(3)  => mem_array(3)(253),
      output(4)  => mem_array(4)(253),
      output(5)  => mem_array(5)(253),
      output(6)  => mem_array(6)(253),
      output(7)  => mem_array(7)(253),
      output(8)  => mem_array(8)(253),
      output(9)  => mem_array(9)(253),
      output(10) => mem_array(10)(253),
      output(11) => mem_array(11)(253),
      output(12) => mem_array(12)(253),
      output(13) => mem_array(13)(253),
      output(14) => mem_array(14)(253),
      output(15) => mem_array(15)(253),
      output(16) => mem_array(16)(253),
      output(17) => mem_array(17)(253),
      output(18) => mem_array(18)(253),
      output(19) => mem_array(19)(253),
      output(20) => mem_array(20)(253),
      output(21) => mem_array(21)(253),
      output(22) => mem_array(22)(253),
      output(23) => mem_array(23)(253),
      output(24) => mem_array(24)(253),
      output(25) => mem_array(25)(253),
      output(26) => mem_array(26)(253),
      output(27) => mem_array(27)(253),
      output(28) => mem_array(28)(253),
      output(29) => mem_array(29)(253),
      output(30) => mem_array(30)(253),
      output(31) => mem_array(31)(253),
      output(32) => mem_array(32)(253),
      output(33) => mem_array(33)(253),
      output(34) => mem_array(34)(253),
      output(35) => mem_array(35)(253)
      );
  rom254 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(254),
      output(0)  => mem_array(0)(254),
      output(1)  => mem_array(1)(254),
      output(2)  => mem_array(2)(254),
      output(3)  => mem_array(3)(254),
      output(4)  => mem_array(4)(254),
      output(5)  => mem_array(5)(254),
      output(6)  => mem_array(6)(254),
      output(7)  => mem_array(7)(254),
      output(8)  => mem_array(8)(254),
      output(9)  => mem_array(9)(254),
      output(10) => mem_array(10)(254),
      output(11) => mem_array(11)(254),
      output(12) => mem_array(12)(254),
      output(13) => mem_array(13)(254),
      output(14) => mem_array(14)(254),
      output(15) => mem_array(15)(254),
      output(16) => mem_array(16)(254),
      output(17) => mem_array(17)(254),
      output(18) => mem_array(18)(254),
      output(19) => mem_array(19)(254),
      output(20) => mem_array(20)(254),
      output(21) => mem_array(21)(254),
      output(22) => mem_array(22)(254),
      output(23) => mem_array(23)(254),
      output(24) => mem_array(24)(254),
      output(25) => mem_array(25)(254),
      output(26) => mem_array(26)(254),
      output(27) => mem_array(27)(254),
      output(28) => mem_array(28)(254),
      output(29) => mem_array(29)(254),
      output(30) => mem_array(30)(254),
      output(31) => mem_array(31)(254),
      output(32) => mem_array(32)(254),
      output(33) => mem_array(33)(254),
      output(34) => mem_array(34)(254),
      output(35) => mem_array(35)(254)
      );
  rom255 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(255),
      output(0)  => mem_array(0)(255),
      output(1)  => mem_array(1)(255),
      output(2)  => mem_array(2)(255),
      output(3)  => mem_array(3)(255),
      output(4)  => mem_array(4)(255),
      output(5)  => mem_array(5)(255),
      output(6)  => mem_array(6)(255),
      output(7)  => mem_array(7)(255),
      output(8)  => mem_array(8)(255),
      output(9)  => mem_array(9)(255),
      output(10) => mem_array(10)(255),
      output(11) => mem_array(11)(255),
      output(12) => mem_array(12)(255),
      output(13) => mem_array(13)(255),
      output(14) => mem_array(14)(255),
      output(15) => mem_array(15)(255),
      output(16) => mem_array(16)(255),
      output(17) => mem_array(17)(255),
      output(18) => mem_array(18)(255),
      output(19) => mem_array(19)(255),
      output(20) => mem_array(20)(255),
      output(21) => mem_array(21)(255),
      output(22) => mem_array(22)(255),
      output(23) => mem_array(23)(255),
      output(24) => mem_array(24)(255),
      output(25) => mem_array(25)(255),
      output(26) => mem_array(26)(255),
      output(27) => mem_array(27)(255),
      output(28) => mem_array(28)(255),
      output(29) => mem_array(29)(255),
      output(30) => mem_array(30)(255),
      output(31) => mem_array(31)(255),
      output(32) => mem_array(32)(255),
      output(33) => mem_array(33)(255),
      output(34) => mem_array(34)(255),
      output(35) => mem_array(35)(255)
      );
  rom256 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(256),
      output(0)  => mem_array(0)(256),
      output(1)  => mem_array(1)(256),
      output(2)  => mem_array(2)(256),
      output(3)  => mem_array(3)(256),
      output(4)  => mem_array(4)(256),
      output(5)  => mem_array(5)(256),
      output(6)  => mem_array(6)(256),
      output(7)  => mem_array(7)(256),
      output(8)  => mem_array(8)(256),
      output(9)  => mem_array(9)(256),
      output(10) => mem_array(10)(256),
      output(11) => mem_array(11)(256),
      output(12) => mem_array(12)(256),
      output(13) => mem_array(13)(256),
      output(14) => mem_array(14)(256),
      output(15) => mem_array(15)(256),
      output(16) => mem_array(16)(256),
      output(17) => mem_array(17)(256),
      output(18) => mem_array(18)(256),
      output(19) => mem_array(19)(256),
      output(20) => mem_array(20)(256),
      output(21) => mem_array(21)(256),
      output(22) => mem_array(22)(256),
      output(23) => mem_array(23)(256),
      output(24) => mem_array(24)(256),
      output(25) => mem_array(25)(256),
      output(26) => mem_array(26)(256),
      output(27) => mem_array(27)(256),
      output(28) => mem_array(28)(256),
      output(29) => mem_array(29)(256),
      output(30) => mem_array(30)(256),
      output(31) => mem_array(31)(256),
      output(32) => mem_array(32)(256),
      output(33) => mem_array(33)(256),
      output(34) => mem_array(34)(256),
      output(35) => mem_array(35)(256)
      );
  rom257 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(257),
      output(0)  => mem_array(0)(257),
      output(1)  => mem_array(1)(257),
      output(2)  => mem_array(2)(257),
      output(3)  => mem_array(3)(257),
      output(4)  => mem_array(4)(257),
      output(5)  => mem_array(5)(257),
      output(6)  => mem_array(6)(257),
      output(7)  => mem_array(7)(257),
      output(8)  => mem_array(8)(257),
      output(9)  => mem_array(9)(257),
      output(10) => mem_array(10)(257),
      output(11) => mem_array(11)(257),
      output(12) => mem_array(12)(257),
      output(13) => mem_array(13)(257),
      output(14) => mem_array(14)(257),
      output(15) => mem_array(15)(257),
      output(16) => mem_array(16)(257),
      output(17) => mem_array(17)(257),
      output(18) => mem_array(18)(257),
      output(19) => mem_array(19)(257),
      output(20) => mem_array(20)(257),
      output(21) => mem_array(21)(257),
      output(22) => mem_array(22)(257),
      output(23) => mem_array(23)(257),
      output(24) => mem_array(24)(257),
      output(25) => mem_array(25)(257),
      output(26) => mem_array(26)(257),
      output(27) => mem_array(27)(257),
      output(28) => mem_array(28)(257),
      output(29) => mem_array(29)(257),
      output(30) => mem_array(30)(257),
      output(31) => mem_array(31)(257),
      output(32) => mem_array(32)(257),
      output(33) => mem_array(33)(257),
      output(34) => mem_array(34)(257),
      output(35) => mem_array(35)(257)
      );
  rom258 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(258),
      output(0)  => mem_array(0)(258),
      output(1)  => mem_array(1)(258),
      output(2)  => mem_array(2)(258),
      output(3)  => mem_array(3)(258),
      output(4)  => mem_array(4)(258),
      output(5)  => mem_array(5)(258),
      output(6)  => mem_array(6)(258),
      output(7)  => mem_array(7)(258),
      output(8)  => mem_array(8)(258),
      output(9)  => mem_array(9)(258),
      output(10) => mem_array(10)(258),
      output(11) => mem_array(11)(258),
      output(12) => mem_array(12)(258),
      output(13) => mem_array(13)(258),
      output(14) => mem_array(14)(258),
      output(15) => mem_array(15)(258),
      output(16) => mem_array(16)(258),
      output(17) => mem_array(17)(258),
      output(18) => mem_array(18)(258),
      output(19) => mem_array(19)(258),
      output(20) => mem_array(20)(258),
      output(21) => mem_array(21)(258),
      output(22) => mem_array(22)(258),
      output(23) => mem_array(23)(258),
      output(24) => mem_array(24)(258),
      output(25) => mem_array(25)(258),
      output(26) => mem_array(26)(258),
      output(27) => mem_array(27)(258),
      output(28) => mem_array(28)(258),
      output(29) => mem_array(29)(258),
      output(30) => mem_array(30)(258),
      output(31) => mem_array(31)(258),
      output(32) => mem_array(32)(258),
      output(33) => mem_array(33)(258),
      output(34) => mem_array(34)(258),
      output(35) => mem_array(35)(258)
      );
  rom259 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(259),
      output(0)  => mem_array(0)(259),
      output(1)  => mem_array(1)(259),
      output(2)  => mem_array(2)(259),
      output(3)  => mem_array(3)(259),
      output(4)  => mem_array(4)(259),
      output(5)  => mem_array(5)(259),
      output(6)  => mem_array(6)(259),
      output(7)  => mem_array(7)(259),
      output(8)  => mem_array(8)(259),
      output(9)  => mem_array(9)(259),
      output(10) => mem_array(10)(259),
      output(11) => mem_array(11)(259),
      output(12) => mem_array(12)(259),
      output(13) => mem_array(13)(259),
      output(14) => mem_array(14)(259),
      output(15) => mem_array(15)(259),
      output(16) => mem_array(16)(259),
      output(17) => mem_array(17)(259),
      output(18) => mem_array(18)(259),
      output(19) => mem_array(19)(259),
      output(20) => mem_array(20)(259),
      output(21) => mem_array(21)(259),
      output(22) => mem_array(22)(259),
      output(23) => mem_array(23)(259),
      output(24) => mem_array(24)(259),
      output(25) => mem_array(25)(259),
      output(26) => mem_array(26)(259),
      output(27) => mem_array(27)(259),
      output(28) => mem_array(28)(259),
      output(29) => mem_array(29)(259),
      output(30) => mem_array(30)(259),
      output(31) => mem_array(31)(259),
      output(32) => mem_array(32)(259),
      output(33) => mem_array(33)(259),
      output(34) => mem_array(34)(259),
      output(35) => mem_array(35)(259)
      );
  rom260 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(260),
      output(0)  => mem_array(0)(260),
      output(1)  => mem_array(1)(260),
      output(2)  => mem_array(2)(260),
      output(3)  => mem_array(3)(260),
      output(4)  => mem_array(4)(260),
      output(5)  => mem_array(5)(260),
      output(6)  => mem_array(6)(260),
      output(7)  => mem_array(7)(260),
      output(8)  => mem_array(8)(260),
      output(9)  => mem_array(9)(260),
      output(10) => mem_array(10)(260),
      output(11) => mem_array(11)(260),
      output(12) => mem_array(12)(260),
      output(13) => mem_array(13)(260),
      output(14) => mem_array(14)(260),
      output(15) => mem_array(15)(260),
      output(16) => mem_array(16)(260),
      output(17) => mem_array(17)(260),
      output(18) => mem_array(18)(260),
      output(19) => mem_array(19)(260),
      output(20) => mem_array(20)(260),
      output(21) => mem_array(21)(260),
      output(22) => mem_array(22)(260),
      output(23) => mem_array(23)(260),
      output(24) => mem_array(24)(260),
      output(25) => mem_array(25)(260),
      output(26) => mem_array(26)(260),
      output(27) => mem_array(27)(260),
      output(28) => mem_array(28)(260),
      output(29) => mem_array(29)(260),
      output(30) => mem_array(30)(260),
      output(31) => mem_array(31)(260),
      output(32) => mem_array(32)(260),
      output(33) => mem_array(33)(260),
      output(34) => mem_array(34)(260),
      output(35) => mem_array(35)(260)
      );
  rom261 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(261),
      output(0)  => mem_array(0)(261),
      output(1)  => mem_array(1)(261),
      output(2)  => mem_array(2)(261),
      output(3)  => mem_array(3)(261),
      output(4)  => mem_array(4)(261),
      output(5)  => mem_array(5)(261),
      output(6)  => mem_array(6)(261),
      output(7)  => mem_array(7)(261),
      output(8)  => mem_array(8)(261),
      output(9)  => mem_array(9)(261),
      output(10) => mem_array(10)(261),
      output(11) => mem_array(11)(261),
      output(12) => mem_array(12)(261),
      output(13) => mem_array(13)(261),
      output(14) => mem_array(14)(261),
      output(15) => mem_array(15)(261),
      output(16) => mem_array(16)(261),
      output(17) => mem_array(17)(261),
      output(18) => mem_array(18)(261),
      output(19) => mem_array(19)(261),
      output(20) => mem_array(20)(261),
      output(21) => mem_array(21)(261),
      output(22) => mem_array(22)(261),
      output(23) => mem_array(23)(261),
      output(24) => mem_array(24)(261),
      output(25) => mem_array(25)(261),
      output(26) => mem_array(26)(261),
      output(27) => mem_array(27)(261),
      output(28) => mem_array(28)(261),
      output(29) => mem_array(29)(261),
      output(30) => mem_array(30)(261),
      output(31) => mem_array(31)(261),
      output(32) => mem_array(32)(261),
      output(33) => mem_array(33)(261),
      output(34) => mem_array(34)(261),
      output(35) => mem_array(35)(261)
      );
  rom262 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(262),
      output(0)  => mem_array(0)(262),
      output(1)  => mem_array(1)(262),
      output(2)  => mem_array(2)(262),
      output(3)  => mem_array(3)(262),
      output(4)  => mem_array(4)(262),
      output(5)  => mem_array(5)(262),
      output(6)  => mem_array(6)(262),
      output(7)  => mem_array(7)(262),
      output(8)  => mem_array(8)(262),
      output(9)  => mem_array(9)(262),
      output(10) => mem_array(10)(262),
      output(11) => mem_array(11)(262),
      output(12) => mem_array(12)(262),
      output(13) => mem_array(13)(262),
      output(14) => mem_array(14)(262),
      output(15) => mem_array(15)(262),
      output(16) => mem_array(16)(262),
      output(17) => mem_array(17)(262),
      output(18) => mem_array(18)(262),
      output(19) => mem_array(19)(262),
      output(20) => mem_array(20)(262),
      output(21) => mem_array(21)(262),
      output(22) => mem_array(22)(262),
      output(23) => mem_array(23)(262),
      output(24) => mem_array(24)(262),
      output(25) => mem_array(25)(262),
      output(26) => mem_array(26)(262),
      output(27) => mem_array(27)(262),
      output(28) => mem_array(28)(262),
      output(29) => mem_array(29)(262),
      output(30) => mem_array(30)(262),
      output(31) => mem_array(31)(262),
      output(32) => mem_array(32)(262),
      output(33) => mem_array(33)(262),
      output(34) => mem_array(34)(262),
      output(35) => mem_array(35)(262)
      );
  rom263 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(263),
      output(0)  => mem_array(0)(263),
      output(1)  => mem_array(1)(263),
      output(2)  => mem_array(2)(263),
      output(3)  => mem_array(3)(263),
      output(4)  => mem_array(4)(263),
      output(5)  => mem_array(5)(263),
      output(6)  => mem_array(6)(263),
      output(7)  => mem_array(7)(263),
      output(8)  => mem_array(8)(263),
      output(9)  => mem_array(9)(263),
      output(10) => mem_array(10)(263),
      output(11) => mem_array(11)(263),
      output(12) => mem_array(12)(263),
      output(13) => mem_array(13)(263),
      output(14) => mem_array(14)(263),
      output(15) => mem_array(15)(263),
      output(16) => mem_array(16)(263),
      output(17) => mem_array(17)(263),
      output(18) => mem_array(18)(263),
      output(19) => mem_array(19)(263),
      output(20) => mem_array(20)(263),
      output(21) => mem_array(21)(263),
      output(22) => mem_array(22)(263),
      output(23) => mem_array(23)(263),
      output(24) => mem_array(24)(263),
      output(25) => mem_array(25)(263),
      output(26) => mem_array(26)(263),
      output(27) => mem_array(27)(263),
      output(28) => mem_array(28)(263),
      output(29) => mem_array(29)(263),
      output(30) => mem_array(30)(263),
      output(31) => mem_array(31)(263),
      output(32) => mem_array(32)(263),
      output(33) => mem_array(33)(263),
      output(34) => mem_array(34)(263),
      output(35) => mem_array(35)(263)
      );
  rom264 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(264),
      output(0)  => mem_array(0)(264),
      output(1)  => mem_array(1)(264),
      output(2)  => mem_array(2)(264),
      output(3)  => mem_array(3)(264),
      output(4)  => mem_array(4)(264),
      output(5)  => mem_array(5)(264),
      output(6)  => mem_array(6)(264),
      output(7)  => mem_array(7)(264),
      output(8)  => mem_array(8)(264),
      output(9)  => mem_array(9)(264),
      output(10) => mem_array(10)(264),
      output(11) => mem_array(11)(264),
      output(12) => mem_array(12)(264),
      output(13) => mem_array(13)(264),
      output(14) => mem_array(14)(264),
      output(15) => mem_array(15)(264),
      output(16) => mem_array(16)(264),
      output(17) => mem_array(17)(264),
      output(18) => mem_array(18)(264),
      output(19) => mem_array(19)(264),
      output(20) => mem_array(20)(264),
      output(21) => mem_array(21)(264),
      output(22) => mem_array(22)(264),
      output(23) => mem_array(23)(264),
      output(24) => mem_array(24)(264),
      output(25) => mem_array(25)(264),
      output(26) => mem_array(26)(264),
      output(27) => mem_array(27)(264),
      output(28) => mem_array(28)(264),
      output(29) => mem_array(29)(264),
      output(30) => mem_array(30)(264),
      output(31) => mem_array(31)(264),
      output(32) => mem_array(32)(264),
      output(33) => mem_array(33)(264),
      output(34) => mem_array(34)(264),
      output(35) => mem_array(35)(264)
      );
  rom265 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(265),
      output(0)  => mem_array(0)(265),
      output(1)  => mem_array(1)(265),
      output(2)  => mem_array(2)(265),
      output(3)  => mem_array(3)(265),
      output(4)  => mem_array(4)(265),
      output(5)  => mem_array(5)(265),
      output(6)  => mem_array(6)(265),
      output(7)  => mem_array(7)(265),
      output(8)  => mem_array(8)(265),
      output(9)  => mem_array(9)(265),
      output(10) => mem_array(10)(265),
      output(11) => mem_array(11)(265),
      output(12) => mem_array(12)(265),
      output(13) => mem_array(13)(265),
      output(14) => mem_array(14)(265),
      output(15) => mem_array(15)(265),
      output(16) => mem_array(16)(265),
      output(17) => mem_array(17)(265),
      output(18) => mem_array(18)(265),
      output(19) => mem_array(19)(265),
      output(20) => mem_array(20)(265),
      output(21) => mem_array(21)(265),
      output(22) => mem_array(22)(265),
      output(23) => mem_array(23)(265),
      output(24) => mem_array(24)(265),
      output(25) => mem_array(25)(265),
      output(26) => mem_array(26)(265),
      output(27) => mem_array(27)(265),
      output(28) => mem_array(28)(265),
      output(29) => mem_array(29)(265),
      output(30) => mem_array(30)(265),
      output(31) => mem_array(31)(265),
      output(32) => mem_array(32)(265),
      output(33) => mem_array(33)(265),
      output(34) => mem_array(34)(265),
      output(35) => mem_array(35)(265)
      );
  rom266 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(266),
      output(0)  => mem_array(0)(266),
      output(1)  => mem_array(1)(266),
      output(2)  => mem_array(2)(266),
      output(3)  => mem_array(3)(266),
      output(4)  => mem_array(4)(266),
      output(5)  => mem_array(5)(266),
      output(6)  => mem_array(6)(266),
      output(7)  => mem_array(7)(266),
      output(8)  => mem_array(8)(266),
      output(9)  => mem_array(9)(266),
      output(10) => mem_array(10)(266),
      output(11) => mem_array(11)(266),
      output(12) => mem_array(12)(266),
      output(13) => mem_array(13)(266),
      output(14) => mem_array(14)(266),
      output(15) => mem_array(15)(266),
      output(16) => mem_array(16)(266),
      output(17) => mem_array(17)(266),
      output(18) => mem_array(18)(266),
      output(19) => mem_array(19)(266),
      output(20) => mem_array(20)(266),
      output(21) => mem_array(21)(266),
      output(22) => mem_array(22)(266),
      output(23) => mem_array(23)(266),
      output(24) => mem_array(24)(266),
      output(25) => mem_array(25)(266),
      output(26) => mem_array(26)(266),
      output(27) => mem_array(27)(266),
      output(28) => mem_array(28)(266),
      output(29) => mem_array(29)(266),
      output(30) => mem_array(30)(266),
      output(31) => mem_array(31)(266),
      output(32) => mem_array(32)(266),
      output(33) => mem_array(33)(266),
      output(34) => mem_array(34)(266),
      output(35) => mem_array(35)(266)
      );
  rom267 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(267),
      output(0)  => mem_array(0)(267),
      output(1)  => mem_array(1)(267),
      output(2)  => mem_array(2)(267),
      output(3)  => mem_array(3)(267),
      output(4)  => mem_array(4)(267),
      output(5)  => mem_array(5)(267),
      output(6)  => mem_array(6)(267),
      output(7)  => mem_array(7)(267),
      output(8)  => mem_array(8)(267),
      output(9)  => mem_array(9)(267),
      output(10) => mem_array(10)(267),
      output(11) => mem_array(11)(267),
      output(12) => mem_array(12)(267),
      output(13) => mem_array(13)(267),
      output(14) => mem_array(14)(267),
      output(15) => mem_array(15)(267),
      output(16) => mem_array(16)(267),
      output(17) => mem_array(17)(267),
      output(18) => mem_array(18)(267),
      output(19) => mem_array(19)(267),
      output(20) => mem_array(20)(267),
      output(21) => mem_array(21)(267),
      output(22) => mem_array(22)(267),
      output(23) => mem_array(23)(267),
      output(24) => mem_array(24)(267),
      output(25) => mem_array(25)(267),
      output(26) => mem_array(26)(267),
      output(27) => mem_array(27)(267),
      output(28) => mem_array(28)(267),
      output(29) => mem_array(29)(267),
      output(30) => mem_array(30)(267),
      output(31) => mem_array(31)(267),
      output(32) => mem_array(32)(267),
      output(33) => mem_array(33)(267),
      output(34) => mem_array(34)(267),
      output(35) => mem_array(35)(267)
      );
  rom268 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(268),
      output(0)  => mem_array(0)(268),
      output(1)  => mem_array(1)(268),
      output(2)  => mem_array(2)(268),
      output(3)  => mem_array(3)(268),
      output(4)  => mem_array(4)(268),
      output(5)  => mem_array(5)(268),
      output(6)  => mem_array(6)(268),
      output(7)  => mem_array(7)(268),
      output(8)  => mem_array(8)(268),
      output(9)  => mem_array(9)(268),
      output(10) => mem_array(10)(268),
      output(11) => mem_array(11)(268),
      output(12) => mem_array(12)(268),
      output(13) => mem_array(13)(268),
      output(14) => mem_array(14)(268),
      output(15) => mem_array(15)(268),
      output(16) => mem_array(16)(268),
      output(17) => mem_array(17)(268),
      output(18) => mem_array(18)(268),
      output(19) => mem_array(19)(268),
      output(20) => mem_array(20)(268),
      output(21) => mem_array(21)(268),
      output(22) => mem_array(22)(268),
      output(23) => mem_array(23)(268),
      output(24) => mem_array(24)(268),
      output(25) => mem_array(25)(268),
      output(26) => mem_array(26)(268),
      output(27) => mem_array(27)(268),
      output(28) => mem_array(28)(268),
      output(29) => mem_array(29)(268),
      output(30) => mem_array(30)(268),
      output(31) => mem_array(31)(268),
      output(32) => mem_array(32)(268),
      output(33) => mem_array(33)(268),
      output(34) => mem_array(34)(268),
      output(35) => mem_array(35)(268)
      );
  rom269 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(269),
      output(0)  => mem_array(0)(269),
      output(1)  => mem_array(1)(269),
      output(2)  => mem_array(2)(269),
      output(3)  => mem_array(3)(269),
      output(4)  => mem_array(4)(269),
      output(5)  => mem_array(5)(269),
      output(6)  => mem_array(6)(269),
      output(7)  => mem_array(7)(269),
      output(8)  => mem_array(8)(269),
      output(9)  => mem_array(9)(269),
      output(10) => mem_array(10)(269),
      output(11) => mem_array(11)(269),
      output(12) => mem_array(12)(269),
      output(13) => mem_array(13)(269),
      output(14) => mem_array(14)(269),
      output(15) => mem_array(15)(269),
      output(16) => mem_array(16)(269),
      output(17) => mem_array(17)(269),
      output(18) => mem_array(18)(269),
      output(19) => mem_array(19)(269),
      output(20) => mem_array(20)(269),
      output(21) => mem_array(21)(269),
      output(22) => mem_array(22)(269),
      output(23) => mem_array(23)(269),
      output(24) => mem_array(24)(269),
      output(25) => mem_array(25)(269),
      output(26) => mem_array(26)(269),
      output(27) => mem_array(27)(269),
      output(28) => mem_array(28)(269),
      output(29) => mem_array(29)(269),
      output(30) => mem_array(30)(269),
      output(31) => mem_array(31)(269),
      output(32) => mem_array(32)(269),
      output(33) => mem_array(33)(269),
      output(34) => mem_array(34)(269),
      output(35) => mem_array(35)(269)
      );
  rom270 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(270),
      output(0)  => mem_array(0)(270),
      output(1)  => mem_array(1)(270),
      output(2)  => mem_array(2)(270),
      output(3)  => mem_array(3)(270),
      output(4)  => mem_array(4)(270),
      output(5)  => mem_array(5)(270),
      output(6)  => mem_array(6)(270),
      output(7)  => mem_array(7)(270),
      output(8)  => mem_array(8)(270),
      output(9)  => mem_array(9)(270),
      output(10) => mem_array(10)(270),
      output(11) => mem_array(11)(270),
      output(12) => mem_array(12)(270),
      output(13) => mem_array(13)(270),
      output(14) => mem_array(14)(270),
      output(15) => mem_array(15)(270),
      output(16) => mem_array(16)(270),
      output(17) => mem_array(17)(270),
      output(18) => mem_array(18)(270),
      output(19) => mem_array(19)(270),
      output(20) => mem_array(20)(270),
      output(21) => mem_array(21)(270),
      output(22) => mem_array(22)(270),
      output(23) => mem_array(23)(270),
      output(24) => mem_array(24)(270),
      output(25) => mem_array(25)(270),
      output(26) => mem_array(26)(270),
      output(27) => mem_array(27)(270),
      output(28) => mem_array(28)(270),
      output(29) => mem_array(29)(270),
      output(30) => mem_array(30)(270),
      output(31) => mem_array(31)(270),
      output(32) => mem_array(32)(270),
      output(33) => mem_array(33)(270),
      output(34) => mem_array(34)(270),
      output(35) => mem_array(35)(270)
      );
  rom271 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(271),
      output(0)  => mem_array(0)(271),
      output(1)  => mem_array(1)(271),
      output(2)  => mem_array(2)(271),
      output(3)  => mem_array(3)(271),
      output(4)  => mem_array(4)(271),
      output(5)  => mem_array(5)(271),
      output(6)  => mem_array(6)(271),
      output(7)  => mem_array(7)(271),
      output(8)  => mem_array(8)(271),
      output(9)  => mem_array(9)(271),
      output(10) => mem_array(10)(271),
      output(11) => mem_array(11)(271),
      output(12) => mem_array(12)(271),
      output(13) => mem_array(13)(271),
      output(14) => mem_array(14)(271),
      output(15) => mem_array(15)(271),
      output(16) => mem_array(16)(271),
      output(17) => mem_array(17)(271),
      output(18) => mem_array(18)(271),
      output(19) => mem_array(19)(271),
      output(20) => mem_array(20)(271),
      output(21) => mem_array(21)(271),
      output(22) => mem_array(22)(271),
      output(23) => mem_array(23)(271),
      output(24) => mem_array(24)(271),
      output(25) => mem_array(25)(271),
      output(26) => mem_array(26)(271),
      output(27) => mem_array(27)(271),
      output(28) => mem_array(28)(271),
      output(29) => mem_array(29)(271),
      output(30) => mem_array(30)(271),
      output(31) => mem_array(31)(271),
      output(32) => mem_array(32)(271),
      output(33) => mem_array(33)(271),
      output(34) => mem_array(34)(271),
      output(35) => mem_array(35)(271)
      );
  rom272 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(272),
      output(0)  => mem_array(0)(272),
      output(1)  => mem_array(1)(272),
      output(2)  => mem_array(2)(272),
      output(3)  => mem_array(3)(272),
      output(4)  => mem_array(4)(272),
      output(5)  => mem_array(5)(272),
      output(6)  => mem_array(6)(272),
      output(7)  => mem_array(7)(272),
      output(8)  => mem_array(8)(272),
      output(9)  => mem_array(9)(272),
      output(10) => mem_array(10)(272),
      output(11) => mem_array(11)(272),
      output(12) => mem_array(12)(272),
      output(13) => mem_array(13)(272),
      output(14) => mem_array(14)(272),
      output(15) => mem_array(15)(272),
      output(16) => mem_array(16)(272),
      output(17) => mem_array(17)(272),
      output(18) => mem_array(18)(272),
      output(19) => mem_array(19)(272),
      output(20) => mem_array(20)(272),
      output(21) => mem_array(21)(272),
      output(22) => mem_array(22)(272),
      output(23) => mem_array(23)(272),
      output(24) => mem_array(24)(272),
      output(25) => mem_array(25)(272),
      output(26) => mem_array(26)(272),
      output(27) => mem_array(27)(272),
      output(28) => mem_array(28)(272),
      output(29) => mem_array(29)(272),
      output(30) => mem_array(30)(272),
      output(31) => mem_array(31)(272),
      output(32) => mem_array(32)(272),
      output(33) => mem_array(33)(272),
      output(34) => mem_array(34)(272),
      output(35) => mem_array(35)(272)
      );
  rom273 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(273),
      output(0)  => mem_array(0)(273),
      output(1)  => mem_array(1)(273),
      output(2)  => mem_array(2)(273),
      output(3)  => mem_array(3)(273),
      output(4)  => mem_array(4)(273),
      output(5)  => mem_array(5)(273),
      output(6)  => mem_array(6)(273),
      output(7)  => mem_array(7)(273),
      output(8)  => mem_array(8)(273),
      output(9)  => mem_array(9)(273),
      output(10) => mem_array(10)(273),
      output(11) => mem_array(11)(273),
      output(12) => mem_array(12)(273),
      output(13) => mem_array(13)(273),
      output(14) => mem_array(14)(273),
      output(15) => mem_array(15)(273),
      output(16) => mem_array(16)(273),
      output(17) => mem_array(17)(273),
      output(18) => mem_array(18)(273),
      output(19) => mem_array(19)(273),
      output(20) => mem_array(20)(273),
      output(21) => mem_array(21)(273),
      output(22) => mem_array(22)(273),
      output(23) => mem_array(23)(273),
      output(24) => mem_array(24)(273),
      output(25) => mem_array(25)(273),
      output(26) => mem_array(26)(273),
      output(27) => mem_array(27)(273),
      output(28) => mem_array(28)(273),
      output(29) => mem_array(29)(273),
      output(30) => mem_array(30)(273),
      output(31) => mem_array(31)(273),
      output(32) => mem_array(32)(273),
      output(33) => mem_array(33)(273),
      output(34) => mem_array(34)(273),
      output(35) => mem_array(35)(273)
      );
  rom274 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(274),
      output(0)  => mem_array(0)(274),
      output(1)  => mem_array(1)(274),
      output(2)  => mem_array(2)(274),
      output(3)  => mem_array(3)(274),
      output(4)  => mem_array(4)(274),
      output(5)  => mem_array(5)(274),
      output(6)  => mem_array(6)(274),
      output(7)  => mem_array(7)(274),
      output(8)  => mem_array(8)(274),
      output(9)  => mem_array(9)(274),
      output(10) => mem_array(10)(274),
      output(11) => mem_array(11)(274),
      output(12) => mem_array(12)(274),
      output(13) => mem_array(13)(274),
      output(14) => mem_array(14)(274),
      output(15) => mem_array(15)(274),
      output(16) => mem_array(16)(274),
      output(17) => mem_array(17)(274),
      output(18) => mem_array(18)(274),
      output(19) => mem_array(19)(274),
      output(20) => mem_array(20)(274),
      output(21) => mem_array(21)(274),
      output(22) => mem_array(22)(274),
      output(23) => mem_array(23)(274),
      output(24) => mem_array(24)(274),
      output(25) => mem_array(25)(274),
      output(26) => mem_array(26)(274),
      output(27) => mem_array(27)(274),
      output(28) => mem_array(28)(274),
      output(29) => mem_array(29)(274),
      output(30) => mem_array(30)(274),
      output(31) => mem_array(31)(274),
      output(32) => mem_array(32)(274),
      output(33) => mem_array(33)(274),
      output(34) => mem_array(34)(274),
      output(35) => mem_array(35)(274)
      );
  rom275 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(275),
      output(0)  => mem_array(0)(275),
      output(1)  => mem_array(1)(275),
      output(2)  => mem_array(2)(275),
      output(3)  => mem_array(3)(275),
      output(4)  => mem_array(4)(275),
      output(5)  => mem_array(5)(275),
      output(6)  => mem_array(6)(275),
      output(7)  => mem_array(7)(275),
      output(8)  => mem_array(8)(275),
      output(9)  => mem_array(9)(275),
      output(10) => mem_array(10)(275),
      output(11) => mem_array(11)(275),
      output(12) => mem_array(12)(275),
      output(13) => mem_array(13)(275),
      output(14) => mem_array(14)(275),
      output(15) => mem_array(15)(275),
      output(16) => mem_array(16)(275),
      output(17) => mem_array(17)(275),
      output(18) => mem_array(18)(275),
      output(19) => mem_array(19)(275),
      output(20) => mem_array(20)(275),
      output(21) => mem_array(21)(275),
      output(22) => mem_array(22)(275),
      output(23) => mem_array(23)(275),
      output(24) => mem_array(24)(275),
      output(25) => mem_array(25)(275),
      output(26) => mem_array(26)(275),
      output(27) => mem_array(27)(275),
      output(28) => mem_array(28)(275),
      output(29) => mem_array(29)(275),
      output(30) => mem_array(30)(275),
      output(31) => mem_array(31)(275),
      output(32) => mem_array(32)(275),
      output(33) => mem_array(33)(275),
      output(34) => mem_array(34)(275),
      output(35) => mem_array(35)(275)
      );
  rom276 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(276),
      output(0)  => mem_array(0)(276),
      output(1)  => mem_array(1)(276),
      output(2)  => mem_array(2)(276),
      output(3)  => mem_array(3)(276),
      output(4)  => mem_array(4)(276),
      output(5)  => mem_array(5)(276),
      output(6)  => mem_array(6)(276),
      output(7)  => mem_array(7)(276),
      output(8)  => mem_array(8)(276),
      output(9)  => mem_array(9)(276),
      output(10) => mem_array(10)(276),
      output(11) => mem_array(11)(276),
      output(12) => mem_array(12)(276),
      output(13) => mem_array(13)(276),
      output(14) => mem_array(14)(276),
      output(15) => mem_array(15)(276),
      output(16) => mem_array(16)(276),
      output(17) => mem_array(17)(276),
      output(18) => mem_array(18)(276),
      output(19) => mem_array(19)(276),
      output(20) => mem_array(20)(276),
      output(21) => mem_array(21)(276),
      output(22) => mem_array(22)(276),
      output(23) => mem_array(23)(276),
      output(24) => mem_array(24)(276),
      output(25) => mem_array(25)(276),
      output(26) => mem_array(26)(276),
      output(27) => mem_array(27)(276),
      output(28) => mem_array(28)(276),
      output(29) => mem_array(29)(276),
      output(30) => mem_array(30)(276),
      output(31) => mem_array(31)(276),
      output(32) => mem_array(32)(276),
      output(33) => mem_array(33)(276),
      output(34) => mem_array(34)(276),
      output(35) => mem_array(35)(276)
      );
  rom277 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(277),
      output(0)  => mem_array(0)(277),
      output(1)  => mem_array(1)(277),
      output(2)  => mem_array(2)(277),
      output(3)  => mem_array(3)(277),
      output(4)  => mem_array(4)(277),
      output(5)  => mem_array(5)(277),
      output(6)  => mem_array(6)(277),
      output(7)  => mem_array(7)(277),
      output(8)  => mem_array(8)(277),
      output(9)  => mem_array(9)(277),
      output(10) => mem_array(10)(277),
      output(11) => mem_array(11)(277),
      output(12) => mem_array(12)(277),
      output(13) => mem_array(13)(277),
      output(14) => mem_array(14)(277),
      output(15) => mem_array(15)(277),
      output(16) => mem_array(16)(277),
      output(17) => mem_array(17)(277),
      output(18) => mem_array(18)(277),
      output(19) => mem_array(19)(277),
      output(20) => mem_array(20)(277),
      output(21) => mem_array(21)(277),
      output(22) => mem_array(22)(277),
      output(23) => mem_array(23)(277),
      output(24) => mem_array(24)(277),
      output(25) => mem_array(25)(277),
      output(26) => mem_array(26)(277),
      output(27) => mem_array(27)(277),
      output(28) => mem_array(28)(277),
      output(29) => mem_array(29)(277),
      output(30) => mem_array(30)(277),
      output(31) => mem_array(31)(277),
      output(32) => mem_array(32)(277),
      output(33) => mem_array(33)(277),
      output(34) => mem_array(34)(277),
      output(35) => mem_array(35)(277)
      );
  rom278 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(278),
      output(0)  => mem_array(0)(278),
      output(1)  => mem_array(1)(278),
      output(2)  => mem_array(2)(278),
      output(3)  => mem_array(3)(278),
      output(4)  => mem_array(4)(278),
      output(5)  => mem_array(5)(278),
      output(6)  => mem_array(6)(278),
      output(7)  => mem_array(7)(278),
      output(8)  => mem_array(8)(278),
      output(9)  => mem_array(9)(278),
      output(10) => mem_array(10)(278),
      output(11) => mem_array(11)(278),
      output(12) => mem_array(12)(278),
      output(13) => mem_array(13)(278),
      output(14) => mem_array(14)(278),
      output(15) => mem_array(15)(278),
      output(16) => mem_array(16)(278),
      output(17) => mem_array(17)(278),
      output(18) => mem_array(18)(278),
      output(19) => mem_array(19)(278),
      output(20) => mem_array(20)(278),
      output(21) => mem_array(21)(278),
      output(22) => mem_array(22)(278),
      output(23) => mem_array(23)(278),
      output(24) => mem_array(24)(278),
      output(25) => mem_array(25)(278),
      output(26) => mem_array(26)(278),
      output(27) => mem_array(27)(278),
      output(28) => mem_array(28)(278),
      output(29) => mem_array(29)(278),
      output(30) => mem_array(30)(278),
      output(31) => mem_array(31)(278),
      output(32) => mem_array(32)(278),
      output(33) => mem_array(33)(278),
      output(34) => mem_array(34)(278),
      output(35) => mem_array(35)(278)
      );
  rom279 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(279),
      output(0)  => mem_array(0)(279),
      output(1)  => mem_array(1)(279),
      output(2)  => mem_array(2)(279),
      output(3)  => mem_array(3)(279),
      output(4)  => mem_array(4)(279),
      output(5)  => mem_array(5)(279),
      output(6)  => mem_array(6)(279),
      output(7)  => mem_array(7)(279),
      output(8)  => mem_array(8)(279),
      output(9)  => mem_array(9)(279),
      output(10) => mem_array(10)(279),
      output(11) => mem_array(11)(279),
      output(12) => mem_array(12)(279),
      output(13) => mem_array(13)(279),
      output(14) => mem_array(14)(279),
      output(15) => mem_array(15)(279),
      output(16) => mem_array(16)(279),
      output(17) => mem_array(17)(279),
      output(18) => mem_array(18)(279),
      output(19) => mem_array(19)(279),
      output(20) => mem_array(20)(279),
      output(21) => mem_array(21)(279),
      output(22) => mem_array(22)(279),
      output(23) => mem_array(23)(279),
      output(24) => mem_array(24)(279),
      output(25) => mem_array(25)(279),
      output(26) => mem_array(26)(279),
      output(27) => mem_array(27)(279),
      output(28) => mem_array(28)(279),
      output(29) => mem_array(29)(279),
      output(30) => mem_array(30)(279),
      output(31) => mem_array(31)(279),
      output(32) => mem_array(32)(279),
      output(33) => mem_array(33)(279),
      output(34) => mem_array(34)(279),
      output(35) => mem_array(35)(279)
      );
  rom280 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000100")
    port map (
      enable_o   => mem_enable_lines(280),
      output(0)  => mem_array(0)(280),
      output(1)  => mem_array(1)(280),
      output(2)  => mem_array(2)(280),
      output(3)  => mem_array(3)(280),
      output(4)  => mem_array(4)(280),
      output(5)  => mem_array(5)(280),
      output(6)  => mem_array(6)(280),
      output(7)  => mem_array(7)(280),
      output(8)  => mem_array(8)(280),
      output(9)  => mem_array(9)(280),
      output(10) => mem_array(10)(280),
      output(11) => mem_array(11)(280),
      output(12) => mem_array(12)(280),
      output(13) => mem_array(13)(280),
      output(14) => mem_array(14)(280),
      output(15) => mem_array(15)(280),
      output(16) => mem_array(16)(280),
      output(17) => mem_array(17)(280),
      output(18) => mem_array(18)(280),
      output(19) => mem_array(19)(280),
      output(20) => mem_array(20)(280),
      output(21) => mem_array(21)(280),
      output(22) => mem_array(22)(280),
      output(23) => mem_array(23)(280),
      output(24) => mem_array(24)(280),
      output(25) => mem_array(25)(280),
      output(26) => mem_array(26)(280),
      output(27) => mem_array(27)(280),
      output(28) => mem_array(28)(280),
      output(29) => mem_array(29)(280),
      output(30) => mem_array(30)(280),
      output(31) => mem_array(31)(280),
      output(32) => mem_array(32)(280),
      output(33) => mem_array(33)(280),
      output(34) => mem_array(34)(280),
      output(35) => mem_array(35)(280)
      );
  rom281 : entity work.rom
    generic map (
      bits  => 36,
      value => "011010000001001011000000000000000000")
    port map (
      enable_o   => mem_enable_lines(281),
      output(0)  => mem_array(0)(281),
      output(1)  => mem_array(1)(281),
      output(2)  => mem_array(2)(281),
      output(3)  => mem_array(3)(281),
      output(4)  => mem_array(4)(281),
      output(5)  => mem_array(5)(281),
      output(6)  => mem_array(6)(281),
      output(7)  => mem_array(7)(281),
      output(8)  => mem_array(8)(281),
      output(9)  => mem_array(9)(281),
      output(10) => mem_array(10)(281),
      output(11) => mem_array(11)(281),
      output(12) => mem_array(12)(281),
      output(13) => mem_array(13)(281),
      output(14) => mem_array(14)(281),
      output(15) => mem_array(15)(281),
      output(16) => mem_array(16)(281),
      output(17) => mem_array(17)(281),
      output(18) => mem_array(18)(281),
      output(19) => mem_array(19)(281),
      output(20) => mem_array(20)(281),
      output(21) => mem_array(21)(281),
      output(22) => mem_array(22)(281),
      output(23) => mem_array(23)(281),
      output(24) => mem_array(24)(281),
      output(25) => mem_array(25)(281),
      output(26) => mem_array(26)(281),
      output(27) => mem_array(27)(281),
      output(28) => mem_array(28)(281),
      output(29) => mem_array(29)(281),
      output(30) => mem_array(30)(281),
      output(31) => mem_array(31)(281),
      output(32) => mem_array(32)(281),
      output(33) => mem_array(33)(281),
      output(34) => mem_array(34)(281),
      output(35) => mem_array(35)(281)
      );
  rom282 : entity work.rom
    generic map (
      bits  => 36,
      value => "010000110000000100101100000000000000")
    port map (
      enable_o   => mem_enable_lines(282),
      output(0)  => mem_array(0)(282),
      output(1)  => mem_array(1)(282),
      output(2)  => mem_array(2)(282),
      output(3)  => mem_array(3)(282),
      output(4)  => mem_array(4)(282),
      output(5)  => mem_array(5)(282),
      output(6)  => mem_array(6)(282),
      output(7)  => mem_array(7)(282),
      output(8)  => mem_array(8)(282),
      output(9)  => mem_array(9)(282),
      output(10) => mem_array(10)(282),
      output(11) => mem_array(11)(282),
      output(12) => mem_array(12)(282),
      output(13) => mem_array(13)(282),
      output(14) => mem_array(14)(282),
      output(15) => mem_array(15)(282),
      output(16) => mem_array(16)(282),
      output(17) => mem_array(17)(282),
      output(18) => mem_array(18)(282),
      output(19) => mem_array(19)(282),
      output(20) => mem_array(20)(282),
      output(21) => mem_array(21)(282),
      output(22) => mem_array(22)(282),
      output(23) => mem_array(23)(282),
      output(24) => mem_array(24)(282),
      output(25) => mem_array(25)(282),
      output(26) => mem_array(26)(282),
      output(27) => mem_array(27)(282),
      output(28) => mem_array(28)(282),
      output(29) => mem_array(29)(282),
      output(30) => mem_array(30)(282),
      output(31) => mem_array(31)(282),
      output(32) => mem_array(32)(282),
      output(33) => mem_array(33)(282),
      output(34) => mem_array(34)(282),
      output(35) => mem_array(35)(282)
      );
  rom283 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000110001000000010010110000000000")
    port map (
      enable_o   => mem_enable_lines(283),
      output(0)  => mem_array(0)(283),
      output(1)  => mem_array(1)(283),
      output(2)  => mem_array(2)(283),
      output(3)  => mem_array(3)(283),
      output(4)  => mem_array(4)(283),
      output(5)  => mem_array(5)(283),
      output(6)  => mem_array(6)(283),
      output(7)  => mem_array(7)(283),
      output(8)  => mem_array(8)(283),
      output(9)  => mem_array(9)(283),
      output(10) => mem_array(10)(283),
      output(11) => mem_array(11)(283),
      output(12) => mem_array(12)(283),
      output(13) => mem_array(13)(283),
      output(14) => mem_array(14)(283),
      output(15) => mem_array(15)(283),
      output(16) => mem_array(16)(283),
      output(17) => mem_array(17)(283),
      output(18) => mem_array(18)(283),
      output(19) => mem_array(19)(283),
      output(20) => mem_array(20)(283),
      output(21) => mem_array(21)(283),
      output(22) => mem_array(22)(283),
      output(23) => mem_array(23)(283),
      output(24) => mem_array(24)(283),
      output(25) => mem_array(25)(283),
      output(26) => mem_array(26)(283),
      output(27) => mem_array(27)(283),
      output(28) => mem_array(28)(283),
      output(29) => mem_array(29)(283),
      output(30) => mem_array(30)(283),
      output(31) => mem_array(31)(283),
      output(32) => mem_array(32)(283),
      output(33) => mem_array(33)(283),
      output(34) => mem_array(34)(283),
      output(35) => mem_array(35)(283)
      );
  rom284 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111110000000000000000000")
    port map (
      enable_o   => mem_enable_lines(284),
      output(0)  => mem_array(0)(284),
      output(1)  => mem_array(1)(284),
      output(2)  => mem_array(2)(284),
      output(3)  => mem_array(3)(284),
      output(4)  => mem_array(4)(284),
      output(5)  => mem_array(5)(284),
      output(6)  => mem_array(6)(284),
      output(7)  => mem_array(7)(284),
      output(8)  => mem_array(8)(284),
      output(9)  => mem_array(9)(284),
      output(10) => mem_array(10)(284),
      output(11) => mem_array(11)(284),
      output(12) => mem_array(12)(284),
      output(13) => mem_array(13)(284),
      output(14) => mem_array(14)(284),
      output(15) => mem_array(15)(284),
      output(16) => mem_array(16)(284),
      output(17) => mem_array(17)(284),
      output(18) => mem_array(18)(284),
      output(19) => mem_array(19)(284),
      output(20) => mem_array(20)(284),
      output(21) => mem_array(21)(284),
      output(22) => mem_array(22)(284),
      output(23) => mem_array(23)(284),
      output(24) => mem_array(24)(284),
      output(25) => mem_array(25)(284),
      output(26) => mem_array(26)(284),
      output(27) => mem_array(27)(284),
      output(28) => mem_array(28)(284),
      output(29) => mem_array(29)(284),
      output(30) => mem_array(30)(284),
      output(31) => mem_array(31)(284),
      output(32) => mem_array(32)(284),
      output(33) => mem_array(33)(284),
      output(34) => mem_array(34)(284),
      output(35) => mem_array(35)(284)
      );
  rom285 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(285),
      output(0)  => mem_array(0)(285),
      output(1)  => mem_array(1)(285),
      output(2)  => mem_array(2)(285),
      output(3)  => mem_array(3)(285),
      output(4)  => mem_array(4)(285),
      output(5)  => mem_array(5)(285),
      output(6)  => mem_array(6)(285),
      output(7)  => mem_array(7)(285),
      output(8)  => mem_array(8)(285),
      output(9)  => mem_array(9)(285),
      output(10) => mem_array(10)(285),
      output(11) => mem_array(11)(285),
      output(12) => mem_array(12)(285),
      output(13) => mem_array(13)(285),
      output(14) => mem_array(14)(285),
      output(15) => mem_array(15)(285),
      output(16) => mem_array(16)(285),
      output(17) => mem_array(17)(285),
      output(18) => mem_array(18)(285),
      output(19) => mem_array(19)(285),
      output(20) => mem_array(20)(285),
      output(21) => mem_array(21)(285),
      output(22) => mem_array(22)(285),
      output(23) => mem_array(23)(285),
      output(24) => mem_array(24)(285),
      output(25) => mem_array(25)(285),
      output(26) => mem_array(26)(285),
      output(27) => mem_array(27)(285),
      output(28) => mem_array(28)(285),
      output(29) => mem_array(29)(285),
      output(30) => mem_array(30)(285),
      output(31) => mem_array(31)(285),
      output(32) => mem_array(32)(285),
      output(33) => mem_array(33)(285),
      output(34) => mem_array(34)(285),
      output(35) => mem_array(35)(285)
      );
  rom286 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000010111100000110110")
    port map (
      enable_o   => mem_enable_lines(286),
      output(0)  => mem_array(0)(286),
      output(1)  => mem_array(1)(286),
      output(2)  => mem_array(2)(286),
      output(3)  => mem_array(3)(286),
      output(4)  => mem_array(4)(286),
      output(5)  => mem_array(5)(286),
      output(6)  => mem_array(6)(286),
      output(7)  => mem_array(7)(286),
      output(8)  => mem_array(8)(286),
      output(9)  => mem_array(9)(286),
      output(10) => mem_array(10)(286),
      output(11) => mem_array(11)(286),
      output(12) => mem_array(12)(286),
      output(13) => mem_array(13)(286),
      output(14) => mem_array(14)(286),
      output(15) => mem_array(15)(286),
      output(16) => mem_array(16)(286),
      output(17) => mem_array(17)(286),
      output(18) => mem_array(18)(286),
      output(19) => mem_array(19)(286),
      output(20) => mem_array(20)(286),
      output(21) => mem_array(21)(286),
      output(22) => mem_array(22)(286),
      output(23) => mem_array(23)(286),
      output(24) => mem_array(24)(286),
      output(25) => mem_array(25)(286),
      output(26) => mem_array(26)(286),
      output(27) => mem_array(27)(286),
      output(28) => mem_array(28)(286),
      output(29) => mem_array(29)(286),
      output(30) => mem_array(30)(286),
      output(31) => mem_array(31)(286),
      output(32) => mem_array(32)(286),
      output(33) => mem_array(33)(286),
      output(34) => mem_array(34)(286),
      output(35) => mem_array(35)(286)
      );
  rom287 : entity work.rom
    generic map (
      bits  => 36,
      value => "010000000001000100000111111100000000")
    port map (
      enable_o   => mem_enable_lines(287),
      output(0)  => mem_array(0)(287),
      output(1)  => mem_array(1)(287),
      output(2)  => mem_array(2)(287),
      output(3)  => mem_array(3)(287),
      output(4)  => mem_array(4)(287),
      output(5)  => mem_array(5)(287),
      output(6)  => mem_array(6)(287),
      output(7)  => mem_array(7)(287),
      output(8)  => mem_array(8)(287),
      output(9)  => mem_array(9)(287),
      output(10) => mem_array(10)(287),
      output(11) => mem_array(11)(287),
      output(12) => mem_array(12)(287),
      output(13) => mem_array(13)(287),
      output(14) => mem_array(14)(287),
      output(15) => mem_array(15)(287),
      output(16) => mem_array(16)(287),
      output(17) => mem_array(17)(287),
      output(18) => mem_array(18)(287),
      output(19) => mem_array(19)(287),
      output(20) => mem_array(20)(287),
      output(21) => mem_array(21)(287),
      output(22) => mem_array(22)(287),
      output(23) => mem_array(23)(287),
      output(24) => mem_array(24)(287),
      output(25) => mem_array(25)(287),
      output(26) => mem_array(26)(287),
      output(27) => mem_array(27)(287),
      output(28) => mem_array(28)(287),
      output(29) => mem_array(29)(287),
      output(30) => mem_array(30)(287),
      output(31) => mem_array(31)(287),
      output(32) => mem_array(32)(287),
      output(33) => mem_array(33)(287),
      output(34) => mem_array(34)(287),
      output(35) => mem_array(35)(287)
      );
  rom288 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(288),
      output(0)  => mem_array(0)(288),
      output(1)  => mem_array(1)(288),
      output(2)  => mem_array(2)(288),
      output(3)  => mem_array(3)(288),
      output(4)  => mem_array(4)(288),
      output(5)  => mem_array(5)(288),
      output(6)  => mem_array(6)(288),
      output(7)  => mem_array(7)(288),
      output(8)  => mem_array(8)(288),
      output(9)  => mem_array(9)(288),
      output(10) => mem_array(10)(288),
      output(11) => mem_array(11)(288),
      output(12) => mem_array(12)(288),
      output(13) => mem_array(13)(288),
      output(14) => mem_array(14)(288),
      output(15) => mem_array(15)(288),
      output(16) => mem_array(16)(288),
      output(17) => mem_array(17)(288),
      output(18) => mem_array(18)(288),
      output(19) => mem_array(19)(288),
      output(20) => mem_array(20)(288),
      output(21) => mem_array(21)(288),
      output(22) => mem_array(22)(288),
      output(23) => mem_array(23)(288),
      output(24) => mem_array(24)(288),
      output(25) => mem_array(25)(288),
      output(26) => mem_array(26)(288),
      output(27) => mem_array(27)(288),
      output(28) => mem_array(28)(288),
      output(29) => mem_array(29)(288),
      output(30) => mem_array(30)(288),
      output(31) => mem_array(31)(288),
      output(32) => mem_array(32)(288),
      output(33) => mem_array(33)(288),
      output(34) => mem_array(34)(288),
      output(35) => mem_array(35)(288)
      );
  rom289 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(289),
      output(0)  => mem_array(0)(289),
      output(1)  => mem_array(1)(289),
      output(2)  => mem_array(2)(289),
      output(3)  => mem_array(3)(289),
      output(4)  => mem_array(4)(289),
      output(5)  => mem_array(5)(289),
      output(6)  => mem_array(6)(289),
      output(7)  => mem_array(7)(289),
      output(8)  => mem_array(8)(289),
      output(9)  => mem_array(9)(289),
      output(10) => mem_array(10)(289),
      output(11) => mem_array(11)(289),
      output(12) => mem_array(12)(289),
      output(13) => mem_array(13)(289),
      output(14) => mem_array(14)(289),
      output(15) => mem_array(15)(289),
      output(16) => mem_array(16)(289),
      output(17) => mem_array(17)(289),
      output(18) => mem_array(18)(289),
      output(19) => mem_array(19)(289),
      output(20) => mem_array(20)(289),
      output(21) => mem_array(21)(289),
      output(22) => mem_array(22)(289),
      output(23) => mem_array(23)(289),
      output(24) => mem_array(24)(289),
      output(25) => mem_array(25)(289),
      output(26) => mem_array(26)(289),
      output(27) => mem_array(27)(289),
      output(28) => mem_array(28)(289),
      output(29) => mem_array(29)(289),
      output(30) => mem_array(30)(289),
      output(31) => mem_array(31)(289),
      output(32) => mem_array(32)(289),
      output(33) => mem_array(33)(289),
      output(34) => mem_array(34)(289),
      output(35) => mem_array(35)(289)
      );
  rom290 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(290),
      output(0)  => mem_array(0)(290),
      output(1)  => mem_array(1)(290),
      output(2)  => mem_array(2)(290),
      output(3)  => mem_array(3)(290),
      output(4)  => mem_array(4)(290),
      output(5)  => mem_array(5)(290),
      output(6)  => mem_array(6)(290),
      output(7)  => mem_array(7)(290),
      output(8)  => mem_array(8)(290),
      output(9)  => mem_array(9)(290),
      output(10) => mem_array(10)(290),
      output(11) => mem_array(11)(290),
      output(12) => mem_array(12)(290),
      output(13) => mem_array(13)(290),
      output(14) => mem_array(14)(290),
      output(15) => mem_array(15)(290),
      output(16) => mem_array(16)(290),
      output(17) => mem_array(17)(290),
      output(18) => mem_array(18)(290),
      output(19) => mem_array(19)(290),
      output(20) => mem_array(20)(290),
      output(21) => mem_array(21)(290),
      output(22) => mem_array(22)(290),
      output(23) => mem_array(23)(290),
      output(24) => mem_array(24)(290),
      output(25) => mem_array(25)(290),
      output(26) => mem_array(26)(290),
      output(27) => mem_array(27)(290),
      output(28) => mem_array(28)(290),
      output(29) => mem_array(29)(290),
      output(30) => mem_array(30)(290),
      output(31) => mem_array(31)(290),
      output(32) => mem_array(32)(290),
      output(33) => mem_array(33)(290),
      output(34) => mem_array(34)(290),
      output(35) => mem_array(35)(290)
      );
  rom291 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(291),
      output(0)  => mem_array(0)(291),
      output(1)  => mem_array(1)(291),
      output(2)  => mem_array(2)(291),
      output(3)  => mem_array(3)(291),
      output(4)  => mem_array(4)(291),
      output(5)  => mem_array(5)(291),
      output(6)  => mem_array(6)(291),
      output(7)  => mem_array(7)(291),
      output(8)  => mem_array(8)(291),
      output(9)  => mem_array(9)(291),
      output(10) => mem_array(10)(291),
      output(11) => mem_array(11)(291),
      output(12) => mem_array(12)(291),
      output(13) => mem_array(13)(291),
      output(14) => mem_array(14)(291),
      output(15) => mem_array(15)(291),
      output(16) => mem_array(16)(291),
      output(17) => mem_array(17)(291),
      output(18) => mem_array(18)(291),
      output(19) => mem_array(19)(291),
      output(20) => mem_array(20)(291),
      output(21) => mem_array(21)(291),
      output(22) => mem_array(22)(291),
      output(23) => mem_array(23)(291),
      output(24) => mem_array(24)(291),
      output(25) => mem_array(25)(291),
      output(26) => mem_array(26)(291),
      output(27) => mem_array(27)(291),
      output(28) => mem_array(28)(291),
      output(29) => mem_array(29)(291),
      output(30) => mem_array(30)(291),
      output(31) => mem_array(31)(291),
      output(32) => mem_array(32)(291),
      output(33) => mem_array(33)(291),
      output(34) => mem_array(34)(291),
      output(35) => mem_array(35)(291)
      );
  rom292 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(292),
      output(0)  => mem_array(0)(292),
      output(1)  => mem_array(1)(292),
      output(2)  => mem_array(2)(292),
      output(3)  => mem_array(3)(292),
      output(4)  => mem_array(4)(292),
      output(5)  => mem_array(5)(292),
      output(6)  => mem_array(6)(292),
      output(7)  => mem_array(7)(292),
      output(8)  => mem_array(8)(292),
      output(9)  => mem_array(9)(292),
      output(10) => mem_array(10)(292),
      output(11) => mem_array(11)(292),
      output(12) => mem_array(12)(292),
      output(13) => mem_array(13)(292),
      output(14) => mem_array(14)(292),
      output(15) => mem_array(15)(292),
      output(16) => mem_array(16)(292),
      output(17) => mem_array(17)(292),
      output(18) => mem_array(18)(292),
      output(19) => mem_array(19)(292),
      output(20) => mem_array(20)(292),
      output(21) => mem_array(21)(292),
      output(22) => mem_array(22)(292),
      output(23) => mem_array(23)(292),
      output(24) => mem_array(24)(292),
      output(25) => mem_array(25)(292),
      output(26) => mem_array(26)(292),
      output(27) => mem_array(27)(292),
      output(28) => mem_array(28)(292),
      output(29) => mem_array(29)(292),
      output(30) => mem_array(30)(292),
      output(31) => mem_array(31)(292),
      output(32) => mem_array(32)(292),
      output(33) => mem_array(33)(292),
      output(34) => mem_array(34)(292),
      output(35) => mem_array(35)(292)
      );
  rom293 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(293),
      output(0)  => mem_array(0)(293),
      output(1)  => mem_array(1)(293),
      output(2)  => mem_array(2)(293),
      output(3)  => mem_array(3)(293),
      output(4)  => mem_array(4)(293),
      output(5)  => mem_array(5)(293),
      output(6)  => mem_array(6)(293),
      output(7)  => mem_array(7)(293),
      output(8)  => mem_array(8)(293),
      output(9)  => mem_array(9)(293),
      output(10) => mem_array(10)(293),
      output(11) => mem_array(11)(293),
      output(12) => mem_array(12)(293),
      output(13) => mem_array(13)(293),
      output(14) => mem_array(14)(293),
      output(15) => mem_array(15)(293),
      output(16) => mem_array(16)(293),
      output(17) => mem_array(17)(293),
      output(18) => mem_array(18)(293),
      output(19) => mem_array(19)(293),
      output(20) => mem_array(20)(293),
      output(21) => mem_array(21)(293),
      output(22) => mem_array(22)(293),
      output(23) => mem_array(23)(293),
      output(24) => mem_array(24)(293),
      output(25) => mem_array(25)(293),
      output(26) => mem_array(26)(293),
      output(27) => mem_array(27)(293),
      output(28) => mem_array(28)(293),
      output(29) => mem_array(29)(293),
      output(30) => mem_array(30)(293),
      output(31) => mem_array(31)(293),
      output(32) => mem_array(32)(293),
      output(33) => mem_array(33)(293),
      output(34) => mem_array(34)(293),
      output(35) => mem_array(35)(293)
      );
  rom294 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(294),
      output(0)  => mem_array(0)(294),
      output(1)  => mem_array(1)(294),
      output(2)  => mem_array(2)(294),
      output(3)  => mem_array(3)(294),
      output(4)  => mem_array(4)(294),
      output(5)  => mem_array(5)(294),
      output(6)  => mem_array(6)(294),
      output(7)  => mem_array(7)(294),
      output(8)  => mem_array(8)(294),
      output(9)  => mem_array(9)(294),
      output(10) => mem_array(10)(294),
      output(11) => mem_array(11)(294),
      output(12) => mem_array(12)(294),
      output(13) => mem_array(13)(294),
      output(14) => mem_array(14)(294),
      output(15) => mem_array(15)(294),
      output(16) => mem_array(16)(294),
      output(17) => mem_array(17)(294),
      output(18) => mem_array(18)(294),
      output(19) => mem_array(19)(294),
      output(20) => mem_array(20)(294),
      output(21) => mem_array(21)(294),
      output(22) => mem_array(22)(294),
      output(23) => mem_array(23)(294),
      output(24) => mem_array(24)(294),
      output(25) => mem_array(25)(294),
      output(26) => mem_array(26)(294),
      output(27) => mem_array(27)(294),
      output(28) => mem_array(28)(294),
      output(29) => mem_array(29)(294),
      output(30) => mem_array(30)(294),
      output(31) => mem_array(31)(294),
      output(32) => mem_array(32)(294),
      output(33) => mem_array(33)(294),
      output(34) => mem_array(34)(294),
      output(35) => mem_array(35)(294)
      );
  rom295 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(295),
      output(0)  => mem_array(0)(295),
      output(1)  => mem_array(1)(295),
      output(2)  => mem_array(2)(295),
      output(3)  => mem_array(3)(295),
      output(4)  => mem_array(4)(295),
      output(5)  => mem_array(5)(295),
      output(6)  => mem_array(6)(295),
      output(7)  => mem_array(7)(295),
      output(8)  => mem_array(8)(295),
      output(9)  => mem_array(9)(295),
      output(10) => mem_array(10)(295),
      output(11) => mem_array(11)(295),
      output(12) => mem_array(12)(295),
      output(13) => mem_array(13)(295),
      output(14) => mem_array(14)(295),
      output(15) => mem_array(15)(295),
      output(16) => mem_array(16)(295),
      output(17) => mem_array(17)(295),
      output(18) => mem_array(18)(295),
      output(19) => mem_array(19)(295),
      output(20) => mem_array(20)(295),
      output(21) => mem_array(21)(295),
      output(22) => mem_array(22)(295),
      output(23) => mem_array(23)(295),
      output(24) => mem_array(24)(295),
      output(25) => mem_array(25)(295),
      output(26) => mem_array(26)(295),
      output(27) => mem_array(27)(295),
      output(28) => mem_array(28)(295),
      output(29) => mem_array(29)(295),
      output(30) => mem_array(30)(295),
      output(31) => mem_array(31)(295),
      output(32) => mem_array(32)(295),
      output(33) => mem_array(33)(295),
      output(34) => mem_array(34)(295),
      output(35) => mem_array(35)(295)
      );
  rom296 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(296),
      output(0)  => mem_array(0)(296),
      output(1)  => mem_array(1)(296),
      output(2)  => mem_array(2)(296),
      output(3)  => mem_array(3)(296),
      output(4)  => mem_array(4)(296),
      output(5)  => mem_array(5)(296),
      output(6)  => mem_array(6)(296),
      output(7)  => mem_array(7)(296),
      output(8)  => mem_array(8)(296),
      output(9)  => mem_array(9)(296),
      output(10) => mem_array(10)(296),
      output(11) => mem_array(11)(296),
      output(12) => mem_array(12)(296),
      output(13) => mem_array(13)(296),
      output(14) => mem_array(14)(296),
      output(15) => mem_array(15)(296),
      output(16) => mem_array(16)(296),
      output(17) => mem_array(17)(296),
      output(18) => mem_array(18)(296),
      output(19) => mem_array(19)(296),
      output(20) => mem_array(20)(296),
      output(21) => mem_array(21)(296),
      output(22) => mem_array(22)(296),
      output(23) => mem_array(23)(296),
      output(24) => mem_array(24)(296),
      output(25) => mem_array(25)(296),
      output(26) => mem_array(26)(296),
      output(27) => mem_array(27)(296),
      output(28) => mem_array(28)(296),
      output(29) => mem_array(29)(296),
      output(30) => mem_array(30)(296),
      output(31) => mem_array(31)(296),
      output(32) => mem_array(32)(296),
      output(33) => mem_array(33)(296),
      output(34) => mem_array(34)(296),
      output(35) => mem_array(35)(296)
      );
  rom297 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(297),
      output(0)  => mem_array(0)(297),
      output(1)  => mem_array(1)(297),
      output(2)  => mem_array(2)(297),
      output(3)  => mem_array(3)(297),
      output(4)  => mem_array(4)(297),
      output(5)  => mem_array(5)(297),
      output(6)  => mem_array(6)(297),
      output(7)  => mem_array(7)(297),
      output(8)  => mem_array(8)(297),
      output(9)  => mem_array(9)(297),
      output(10) => mem_array(10)(297),
      output(11) => mem_array(11)(297),
      output(12) => mem_array(12)(297),
      output(13) => mem_array(13)(297),
      output(14) => mem_array(14)(297),
      output(15) => mem_array(15)(297),
      output(16) => mem_array(16)(297),
      output(17) => mem_array(17)(297),
      output(18) => mem_array(18)(297),
      output(19) => mem_array(19)(297),
      output(20) => mem_array(20)(297),
      output(21) => mem_array(21)(297),
      output(22) => mem_array(22)(297),
      output(23) => mem_array(23)(297),
      output(24) => mem_array(24)(297),
      output(25) => mem_array(25)(297),
      output(26) => mem_array(26)(297),
      output(27) => mem_array(27)(297),
      output(28) => mem_array(28)(297),
      output(29) => mem_array(29)(297),
      output(30) => mem_array(30)(297),
      output(31) => mem_array(31)(297),
      output(32) => mem_array(32)(297),
      output(33) => mem_array(33)(297),
      output(34) => mem_array(34)(297),
      output(35) => mem_array(35)(297)
      );
  rom298 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(298),
      output(0)  => mem_array(0)(298),
      output(1)  => mem_array(1)(298),
      output(2)  => mem_array(2)(298),
      output(3)  => mem_array(3)(298),
      output(4)  => mem_array(4)(298),
      output(5)  => mem_array(5)(298),
      output(6)  => mem_array(6)(298),
      output(7)  => mem_array(7)(298),
      output(8)  => mem_array(8)(298),
      output(9)  => mem_array(9)(298),
      output(10) => mem_array(10)(298),
      output(11) => mem_array(11)(298),
      output(12) => mem_array(12)(298),
      output(13) => mem_array(13)(298),
      output(14) => mem_array(14)(298),
      output(15) => mem_array(15)(298),
      output(16) => mem_array(16)(298),
      output(17) => mem_array(17)(298),
      output(18) => mem_array(18)(298),
      output(19) => mem_array(19)(298),
      output(20) => mem_array(20)(298),
      output(21) => mem_array(21)(298),
      output(22) => mem_array(22)(298),
      output(23) => mem_array(23)(298),
      output(24) => mem_array(24)(298),
      output(25) => mem_array(25)(298),
      output(26) => mem_array(26)(298),
      output(27) => mem_array(27)(298),
      output(28) => mem_array(28)(298),
      output(29) => mem_array(29)(298),
      output(30) => mem_array(30)(298),
      output(31) => mem_array(31)(298),
      output(32) => mem_array(32)(298),
      output(33) => mem_array(33)(298),
      output(34) => mem_array(34)(298),
      output(35) => mem_array(35)(298)
      );
  rom299 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(299),
      output(0)  => mem_array(0)(299),
      output(1)  => mem_array(1)(299),
      output(2)  => mem_array(2)(299),
      output(3)  => mem_array(3)(299),
      output(4)  => mem_array(4)(299),
      output(5)  => mem_array(5)(299),
      output(6)  => mem_array(6)(299),
      output(7)  => mem_array(7)(299),
      output(8)  => mem_array(8)(299),
      output(9)  => mem_array(9)(299),
      output(10) => mem_array(10)(299),
      output(11) => mem_array(11)(299),
      output(12) => mem_array(12)(299),
      output(13) => mem_array(13)(299),
      output(14) => mem_array(14)(299),
      output(15) => mem_array(15)(299),
      output(16) => mem_array(16)(299),
      output(17) => mem_array(17)(299),
      output(18) => mem_array(18)(299),
      output(19) => mem_array(19)(299),
      output(20) => mem_array(20)(299),
      output(21) => mem_array(21)(299),
      output(22) => mem_array(22)(299),
      output(23) => mem_array(23)(299),
      output(24) => mem_array(24)(299),
      output(25) => mem_array(25)(299),
      output(26) => mem_array(26)(299),
      output(27) => mem_array(27)(299),
      output(28) => mem_array(28)(299),
      output(29) => mem_array(29)(299),
      output(30) => mem_array(30)(299),
      output(31) => mem_array(31)(299),
      output(32) => mem_array(32)(299),
      output(33) => mem_array(33)(299),
      output(34) => mem_array(34)(299),
      output(35) => mem_array(35)(299)
      );
  rom300 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(300),
      output(0)  => mem_array(0)(300),
      output(1)  => mem_array(1)(300),
      output(2)  => mem_array(2)(300),
      output(3)  => mem_array(3)(300),
      output(4)  => mem_array(4)(300),
      output(5)  => mem_array(5)(300),
      output(6)  => mem_array(6)(300),
      output(7)  => mem_array(7)(300),
      output(8)  => mem_array(8)(300),
      output(9)  => mem_array(9)(300),
      output(10) => mem_array(10)(300),
      output(11) => mem_array(11)(300),
      output(12) => mem_array(12)(300),
      output(13) => mem_array(13)(300),
      output(14) => mem_array(14)(300),
      output(15) => mem_array(15)(300),
      output(16) => mem_array(16)(300),
      output(17) => mem_array(17)(300),
      output(18) => mem_array(18)(300),
      output(19) => mem_array(19)(300),
      output(20) => mem_array(20)(300),
      output(21) => mem_array(21)(300),
      output(22) => mem_array(22)(300),
      output(23) => mem_array(23)(300),
      output(24) => mem_array(24)(300),
      output(25) => mem_array(25)(300),
      output(26) => mem_array(26)(300),
      output(27) => mem_array(27)(300),
      output(28) => mem_array(28)(300),
      output(29) => mem_array(29)(300),
      output(30) => mem_array(30)(300),
      output(31) => mem_array(31)(300),
      output(32) => mem_array(32)(300),
      output(33) => mem_array(33)(300),
      output(34) => mem_array(34)(300),
      output(35) => mem_array(35)(300)
      );
  rom301 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(301),
      output(0)  => mem_array(0)(301),
      output(1)  => mem_array(1)(301),
      output(2)  => mem_array(2)(301),
      output(3)  => mem_array(3)(301),
      output(4)  => mem_array(4)(301),
      output(5)  => mem_array(5)(301),
      output(6)  => mem_array(6)(301),
      output(7)  => mem_array(7)(301),
      output(8)  => mem_array(8)(301),
      output(9)  => mem_array(9)(301),
      output(10) => mem_array(10)(301),
      output(11) => mem_array(11)(301),
      output(12) => mem_array(12)(301),
      output(13) => mem_array(13)(301),
      output(14) => mem_array(14)(301),
      output(15) => mem_array(15)(301),
      output(16) => mem_array(16)(301),
      output(17) => mem_array(17)(301),
      output(18) => mem_array(18)(301),
      output(19) => mem_array(19)(301),
      output(20) => mem_array(20)(301),
      output(21) => mem_array(21)(301),
      output(22) => mem_array(22)(301),
      output(23) => mem_array(23)(301),
      output(24) => mem_array(24)(301),
      output(25) => mem_array(25)(301),
      output(26) => mem_array(26)(301),
      output(27) => mem_array(27)(301),
      output(28) => mem_array(28)(301),
      output(29) => mem_array(29)(301),
      output(30) => mem_array(30)(301),
      output(31) => mem_array(31)(301),
      output(32) => mem_array(32)(301),
      output(33) => mem_array(33)(301),
      output(34) => mem_array(34)(301),
      output(35) => mem_array(35)(301)
      );
  rom302 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(302),
      output(0)  => mem_array(0)(302),
      output(1)  => mem_array(1)(302),
      output(2)  => mem_array(2)(302),
      output(3)  => mem_array(3)(302),
      output(4)  => mem_array(4)(302),
      output(5)  => mem_array(5)(302),
      output(6)  => mem_array(6)(302),
      output(7)  => mem_array(7)(302),
      output(8)  => mem_array(8)(302),
      output(9)  => mem_array(9)(302),
      output(10) => mem_array(10)(302),
      output(11) => mem_array(11)(302),
      output(12) => mem_array(12)(302),
      output(13) => mem_array(13)(302),
      output(14) => mem_array(14)(302),
      output(15) => mem_array(15)(302),
      output(16) => mem_array(16)(302),
      output(17) => mem_array(17)(302),
      output(18) => mem_array(18)(302),
      output(19) => mem_array(19)(302),
      output(20) => mem_array(20)(302),
      output(21) => mem_array(21)(302),
      output(22) => mem_array(22)(302),
      output(23) => mem_array(23)(302),
      output(24) => mem_array(24)(302),
      output(25) => mem_array(25)(302),
      output(26) => mem_array(26)(302),
      output(27) => mem_array(27)(302),
      output(28) => mem_array(28)(302),
      output(29) => mem_array(29)(302),
      output(30) => mem_array(30)(302),
      output(31) => mem_array(31)(302),
      output(32) => mem_array(32)(302),
      output(33) => mem_array(33)(302),
      output(34) => mem_array(34)(302),
      output(35) => mem_array(35)(302)
      );
  rom303 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(303),
      output(0)  => mem_array(0)(303),
      output(1)  => mem_array(1)(303),
      output(2)  => mem_array(2)(303),
      output(3)  => mem_array(3)(303),
      output(4)  => mem_array(4)(303),
      output(5)  => mem_array(5)(303),
      output(6)  => mem_array(6)(303),
      output(7)  => mem_array(7)(303),
      output(8)  => mem_array(8)(303),
      output(9)  => mem_array(9)(303),
      output(10) => mem_array(10)(303),
      output(11) => mem_array(11)(303),
      output(12) => mem_array(12)(303),
      output(13) => mem_array(13)(303),
      output(14) => mem_array(14)(303),
      output(15) => mem_array(15)(303),
      output(16) => mem_array(16)(303),
      output(17) => mem_array(17)(303),
      output(18) => mem_array(18)(303),
      output(19) => mem_array(19)(303),
      output(20) => mem_array(20)(303),
      output(21) => mem_array(21)(303),
      output(22) => mem_array(22)(303),
      output(23) => mem_array(23)(303),
      output(24) => mem_array(24)(303),
      output(25) => mem_array(25)(303),
      output(26) => mem_array(26)(303),
      output(27) => mem_array(27)(303),
      output(28) => mem_array(28)(303),
      output(29) => mem_array(29)(303),
      output(30) => mem_array(30)(303),
      output(31) => mem_array(31)(303),
      output(32) => mem_array(32)(303),
      output(33) => mem_array(33)(303),
      output(34) => mem_array(34)(303),
      output(35) => mem_array(35)(303)
      );
  rom304 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(304),
      output(0)  => mem_array(0)(304),
      output(1)  => mem_array(1)(304),
      output(2)  => mem_array(2)(304),
      output(3)  => mem_array(3)(304),
      output(4)  => mem_array(4)(304),
      output(5)  => mem_array(5)(304),
      output(6)  => mem_array(6)(304),
      output(7)  => mem_array(7)(304),
      output(8)  => mem_array(8)(304),
      output(9)  => mem_array(9)(304),
      output(10) => mem_array(10)(304),
      output(11) => mem_array(11)(304),
      output(12) => mem_array(12)(304),
      output(13) => mem_array(13)(304),
      output(14) => mem_array(14)(304),
      output(15) => mem_array(15)(304),
      output(16) => mem_array(16)(304),
      output(17) => mem_array(17)(304),
      output(18) => mem_array(18)(304),
      output(19) => mem_array(19)(304),
      output(20) => mem_array(20)(304),
      output(21) => mem_array(21)(304),
      output(22) => mem_array(22)(304),
      output(23) => mem_array(23)(304),
      output(24) => mem_array(24)(304),
      output(25) => mem_array(25)(304),
      output(26) => mem_array(26)(304),
      output(27) => mem_array(27)(304),
      output(28) => mem_array(28)(304),
      output(29) => mem_array(29)(304),
      output(30) => mem_array(30)(304),
      output(31) => mem_array(31)(304),
      output(32) => mem_array(32)(304),
      output(33) => mem_array(33)(304),
      output(34) => mem_array(34)(304),
      output(35) => mem_array(35)(304)
      );
  rom305 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(305),
      output(0)  => mem_array(0)(305),
      output(1)  => mem_array(1)(305),
      output(2)  => mem_array(2)(305),
      output(3)  => mem_array(3)(305),
      output(4)  => mem_array(4)(305),
      output(5)  => mem_array(5)(305),
      output(6)  => mem_array(6)(305),
      output(7)  => mem_array(7)(305),
      output(8)  => mem_array(8)(305),
      output(9)  => mem_array(9)(305),
      output(10) => mem_array(10)(305),
      output(11) => mem_array(11)(305),
      output(12) => mem_array(12)(305),
      output(13) => mem_array(13)(305),
      output(14) => mem_array(14)(305),
      output(15) => mem_array(15)(305),
      output(16) => mem_array(16)(305),
      output(17) => mem_array(17)(305),
      output(18) => mem_array(18)(305),
      output(19) => mem_array(19)(305),
      output(20) => mem_array(20)(305),
      output(21) => mem_array(21)(305),
      output(22) => mem_array(22)(305),
      output(23) => mem_array(23)(305),
      output(24) => mem_array(24)(305),
      output(25) => mem_array(25)(305),
      output(26) => mem_array(26)(305),
      output(27) => mem_array(27)(305),
      output(28) => mem_array(28)(305),
      output(29) => mem_array(29)(305),
      output(30) => mem_array(30)(305),
      output(31) => mem_array(31)(305),
      output(32) => mem_array(32)(305),
      output(33) => mem_array(33)(305),
      output(34) => mem_array(34)(305),
      output(35) => mem_array(35)(305)
      );
  rom306 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(306),
      output(0)  => mem_array(0)(306),
      output(1)  => mem_array(1)(306),
      output(2)  => mem_array(2)(306),
      output(3)  => mem_array(3)(306),
      output(4)  => mem_array(4)(306),
      output(5)  => mem_array(5)(306),
      output(6)  => mem_array(6)(306),
      output(7)  => mem_array(7)(306),
      output(8)  => mem_array(8)(306),
      output(9)  => mem_array(9)(306),
      output(10) => mem_array(10)(306),
      output(11) => mem_array(11)(306),
      output(12) => mem_array(12)(306),
      output(13) => mem_array(13)(306),
      output(14) => mem_array(14)(306),
      output(15) => mem_array(15)(306),
      output(16) => mem_array(16)(306),
      output(17) => mem_array(17)(306),
      output(18) => mem_array(18)(306),
      output(19) => mem_array(19)(306),
      output(20) => mem_array(20)(306),
      output(21) => mem_array(21)(306),
      output(22) => mem_array(22)(306),
      output(23) => mem_array(23)(306),
      output(24) => mem_array(24)(306),
      output(25) => mem_array(25)(306),
      output(26) => mem_array(26)(306),
      output(27) => mem_array(27)(306),
      output(28) => mem_array(28)(306),
      output(29) => mem_array(29)(306),
      output(30) => mem_array(30)(306),
      output(31) => mem_array(31)(306),
      output(32) => mem_array(32)(306),
      output(33) => mem_array(33)(306),
      output(34) => mem_array(34)(306),
      output(35) => mem_array(35)(306)
      );
  rom307 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(307),
      output(0)  => mem_array(0)(307),
      output(1)  => mem_array(1)(307),
      output(2)  => mem_array(2)(307),
      output(3)  => mem_array(3)(307),
      output(4)  => mem_array(4)(307),
      output(5)  => mem_array(5)(307),
      output(6)  => mem_array(6)(307),
      output(7)  => mem_array(7)(307),
      output(8)  => mem_array(8)(307),
      output(9)  => mem_array(9)(307),
      output(10) => mem_array(10)(307),
      output(11) => mem_array(11)(307),
      output(12) => mem_array(12)(307),
      output(13) => mem_array(13)(307),
      output(14) => mem_array(14)(307),
      output(15) => mem_array(15)(307),
      output(16) => mem_array(16)(307),
      output(17) => mem_array(17)(307),
      output(18) => mem_array(18)(307),
      output(19) => mem_array(19)(307),
      output(20) => mem_array(20)(307),
      output(21) => mem_array(21)(307),
      output(22) => mem_array(22)(307),
      output(23) => mem_array(23)(307),
      output(24) => mem_array(24)(307),
      output(25) => mem_array(25)(307),
      output(26) => mem_array(26)(307),
      output(27) => mem_array(27)(307),
      output(28) => mem_array(28)(307),
      output(29) => mem_array(29)(307),
      output(30) => mem_array(30)(307),
      output(31) => mem_array(31)(307),
      output(32) => mem_array(32)(307),
      output(33) => mem_array(33)(307),
      output(34) => mem_array(34)(307),
      output(35) => mem_array(35)(307)
      );
  rom308 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000100001000")
    port map (
      enable_o   => mem_enable_lines(308),
      output(0)  => mem_array(0)(308),
      output(1)  => mem_array(1)(308),
      output(2)  => mem_array(2)(308),
      output(3)  => mem_array(3)(308),
      output(4)  => mem_array(4)(308),
      output(5)  => mem_array(5)(308),
      output(6)  => mem_array(6)(308),
      output(7)  => mem_array(7)(308),
      output(8)  => mem_array(8)(308),
      output(9)  => mem_array(9)(308),
      output(10) => mem_array(10)(308),
      output(11) => mem_array(11)(308),
      output(12) => mem_array(12)(308),
      output(13) => mem_array(13)(308),
      output(14) => mem_array(14)(308),
      output(15) => mem_array(15)(308),
      output(16) => mem_array(16)(308),
      output(17) => mem_array(17)(308),
      output(18) => mem_array(18)(308),
      output(19) => mem_array(19)(308),
      output(20) => mem_array(20)(308),
      output(21) => mem_array(21)(308),
      output(22) => mem_array(22)(308),
      output(23) => mem_array(23)(308),
      output(24) => mem_array(24)(308),
      output(25) => mem_array(25)(308),
      output(26) => mem_array(26)(308),
      output(27) => mem_array(27)(308),
      output(28) => mem_array(28)(308),
      output(29) => mem_array(29)(308),
      output(30) => mem_array(30)(308),
      output(31) => mem_array(31)(308),
      output(32) => mem_array(32)(308),
      output(33) => mem_array(33)(308),
      output(34) => mem_array(34)(308),
      output(35) => mem_array(35)(308)
      );
  rom309 : entity work.rom
    generic map (
      bits  => 36,
      value => "001101010000001000010001000001111111")
    port map (
      enable_o   => mem_enable_lines(309),
      output(0)  => mem_array(0)(309),
      output(1)  => mem_array(1)(309),
      output(2)  => mem_array(2)(309),
      output(3)  => mem_array(3)(309),
      output(4)  => mem_array(4)(309),
      output(5)  => mem_array(5)(309),
      output(6)  => mem_array(6)(309),
      output(7)  => mem_array(7)(309),
      output(8)  => mem_array(8)(309),
      output(9)  => mem_array(9)(309),
      output(10) => mem_array(10)(309),
      output(11) => mem_array(11)(309),
      output(12) => mem_array(12)(309),
      output(13) => mem_array(13)(309),
      output(14) => mem_array(14)(309),
      output(15) => mem_array(15)(309),
      output(16) => mem_array(16)(309),
      output(17) => mem_array(17)(309),
      output(18) => mem_array(18)(309),
      output(19) => mem_array(19)(309),
      output(20) => mem_array(20)(309),
      output(21) => mem_array(21)(309),
      output(22) => mem_array(22)(309),
      output(23) => mem_array(23)(309),
      output(24) => mem_array(24)(309),
      output(25) => mem_array(25)(309),
      output(26) => mem_array(26)(309),
      output(27) => mem_array(27)(309),
      output(28) => mem_array(28)(309),
      output(29) => mem_array(29)(309),
      output(30) => mem_array(30)(309),
      output(31) => mem_array(31)(309),
      output(32) => mem_array(32)(309),
      output(33) => mem_array(33)(309),
      output(34) => mem_array(34)(309),
      output(35) => mem_array(35)(309)
      );
  rom310 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(310),
      output(0)  => mem_array(0)(310),
      output(1)  => mem_array(1)(310),
      output(2)  => mem_array(2)(310),
      output(3)  => mem_array(3)(310),
      output(4)  => mem_array(4)(310),
      output(5)  => mem_array(5)(310),
      output(6)  => mem_array(6)(310),
      output(7)  => mem_array(7)(310),
      output(8)  => mem_array(8)(310),
      output(9)  => mem_array(9)(310),
      output(10) => mem_array(10)(310),
      output(11) => mem_array(11)(310),
      output(12) => mem_array(12)(310),
      output(13) => mem_array(13)(310),
      output(14) => mem_array(14)(310),
      output(15) => mem_array(15)(310),
      output(16) => mem_array(16)(310),
      output(17) => mem_array(17)(310),
      output(18) => mem_array(18)(310),
      output(19) => mem_array(19)(310),
      output(20) => mem_array(20)(310),
      output(21) => mem_array(21)(310),
      output(22) => mem_array(22)(310),
      output(23) => mem_array(23)(310),
      output(24) => mem_array(24)(310),
      output(25) => mem_array(25)(310),
      output(26) => mem_array(26)(310),
      output(27) => mem_array(27)(310),
      output(28) => mem_array(28)(310),
      output(29) => mem_array(29)(310),
      output(30) => mem_array(30)(310),
      output(31) => mem_array(31)(310),
      output(32) => mem_array(32)(310),
      output(33) => mem_array(33)(310),
      output(34) => mem_array(34)(310),
      output(35) => mem_array(35)(310)
      );
  rom311 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(311),
      output(0)  => mem_array(0)(311),
      output(1)  => mem_array(1)(311),
      output(2)  => mem_array(2)(311),
      output(3)  => mem_array(3)(311),
      output(4)  => mem_array(4)(311),
      output(5)  => mem_array(5)(311),
      output(6)  => mem_array(6)(311),
      output(7)  => mem_array(7)(311),
      output(8)  => mem_array(8)(311),
      output(9)  => mem_array(9)(311),
      output(10) => mem_array(10)(311),
      output(11) => mem_array(11)(311),
      output(12) => mem_array(12)(311),
      output(13) => mem_array(13)(311),
      output(14) => mem_array(14)(311),
      output(15) => mem_array(15)(311),
      output(16) => mem_array(16)(311),
      output(17) => mem_array(17)(311),
      output(18) => mem_array(18)(311),
      output(19) => mem_array(19)(311),
      output(20) => mem_array(20)(311),
      output(21) => mem_array(21)(311),
      output(22) => mem_array(22)(311),
      output(23) => mem_array(23)(311),
      output(24) => mem_array(24)(311),
      output(25) => mem_array(25)(311),
      output(26) => mem_array(26)(311),
      output(27) => mem_array(27)(311),
      output(28) => mem_array(28)(311),
      output(29) => mem_array(29)(311),
      output(30) => mem_array(30)(311),
      output(31) => mem_array(31)(311),
      output(32) => mem_array(32)(311),
      output(33) => mem_array(33)(311),
      output(34) => mem_array(34)(311),
      output(35) => mem_array(35)(311)
      );
  rom312 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(312),
      output(0)  => mem_array(0)(312),
      output(1)  => mem_array(1)(312),
      output(2)  => mem_array(2)(312),
      output(3)  => mem_array(3)(312),
      output(4)  => mem_array(4)(312),
      output(5)  => mem_array(5)(312),
      output(6)  => mem_array(6)(312),
      output(7)  => mem_array(7)(312),
      output(8)  => mem_array(8)(312),
      output(9)  => mem_array(9)(312),
      output(10) => mem_array(10)(312),
      output(11) => mem_array(11)(312),
      output(12) => mem_array(12)(312),
      output(13) => mem_array(13)(312),
      output(14) => mem_array(14)(312),
      output(15) => mem_array(15)(312),
      output(16) => mem_array(16)(312),
      output(17) => mem_array(17)(312),
      output(18) => mem_array(18)(312),
      output(19) => mem_array(19)(312),
      output(20) => mem_array(20)(312),
      output(21) => mem_array(21)(312),
      output(22) => mem_array(22)(312),
      output(23) => mem_array(23)(312),
      output(24) => mem_array(24)(312),
      output(25) => mem_array(25)(312),
      output(26) => mem_array(26)(312),
      output(27) => mem_array(27)(312),
      output(28) => mem_array(28)(312),
      output(29) => mem_array(29)(312),
      output(30) => mem_array(30)(312),
      output(31) => mem_array(31)(312),
      output(32) => mem_array(32)(312),
      output(33) => mem_array(33)(312),
      output(34) => mem_array(34)(312),
      output(35) => mem_array(35)(312)
      );
  rom313 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(313),
      output(0)  => mem_array(0)(313),
      output(1)  => mem_array(1)(313),
      output(2)  => mem_array(2)(313),
      output(3)  => mem_array(3)(313),
      output(4)  => mem_array(4)(313),
      output(5)  => mem_array(5)(313),
      output(6)  => mem_array(6)(313),
      output(7)  => mem_array(7)(313),
      output(8)  => mem_array(8)(313),
      output(9)  => mem_array(9)(313),
      output(10) => mem_array(10)(313),
      output(11) => mem_array(11)(313),
      output(12) => mem_array(12)(313),
      output(13) => mem_array(13)(313),
      output(14) => mem_array(14)(313),
      output(15) => mem_array(15)(313),
      output(16) => mem_array(16)(313),
      output(17) => mem_array(17)(313),
      output(18) => mem_array(18)(313),
      output(19) => mem_array(19)(313),
      output(20) => mem_array(20)(313),
      output(21) => mem_array(21)(313),
      output(22) => mem_array(22)(313),
      output(23) => mem_array(23)(313),
      output(24) => mem_array(24)(313),
      output(25) => mem_array(25)(313),
      output(26) => mem_array(26)(313),
      output(27) => mem_array(27)(313),
      output(28) => mem_array(28)(313),
      output(29) => mem_array(29)(313),
      output(30) => mem_array(30)(313),
      output(31) => mem_array(31)(313),
      output(32) => mem_array(32)(313),
      output(33) => mem_array(33)(313),
      output(34) => mem_array(34)(313),
      output(35) => mem_array(35)(313)
      );
  rom314 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(314),
      output(0)  => mem_array(0)(314),
      output(1)  => mem_array(1)(314),
      output(2)  => mem_array(2)(314),
      output(3)  => mem_array(3)(314),
      output(4)  => mem_array(4)(314),
      output(5)  => mem_array(5)(314),
      output(6)  => mem_array(6)(314),
      output(7)  => mem_array(7)(314),
      output(8)  => mem_array(8)(314),
      output(9)  => mem_array(9)(314),
      output(10) => mem_array(10)(314),
      output(11) => mem_array(11)(314),
      output(12) => mem_array(12)(314),
      output(13) => mem_array(13)(314),
      output(14) => mem_array(14)(314),
      output(15) => mem_array(15)(314),
      output(16) => mem_array(16)(314),
      output(17) => mem_array(17)(314),
      output(18) => mem_array(18)(314),
      output(19) => mem_array(19)(314),
      output(20) => mem_array(20)(314),
      output(21) => mem_array(21)(314),
      output(22) => mem_array(22)(314),
      output(23) => mem_array(23)(314),
      output(24) => mem_array(24)(314),
      output(25) => mem_array(25)(314),
      output(26) => mem_array(26)(314),
      output(27) => mem_array(27)(314),
      output(28) => mem_array(28)(314),
      output(29) => mem_array(29)(314),
      output(30) => mem_array(30)(314),
      output(31) => mem_array(31)(314),
      output(32) => mem_array(32)(314),
      output(33) => mem_array(33)(314),
      output(34) => mem_array(34)(314),
      output(35) => mem_array(35)(314)
      );
  rom315 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(315),
      output(0)  => mem_array(0)(315),
      output(1)  => mem_array(1)(315),
      output(2)  => mem_array(2)(315),
      output(3)  => mem_array(3)(315),
      output(4)  => mem_array(4)(315),
      output(5)  => mem_array(5)(315),
      output(6)  => mem_array(6)(315),
      output(7)  => mem_array(7)(315),
      output(8)  => mem_array(8)(315),
      output(9)  => mem_array(9)(315),
      output(10) => mem_array(10)(315),
      output(11) => mem_array(11)(315),
      output(12) => mem_array(12)(315),
      output(13) => mem_array(13)(315),
      output(14) => mem_array(14)(315),
      output(15) => mem_array(15)(315),
      output(16) => mem_array(16)(315),
      output(17) => mem_array(17)(315),
      output(18) => mem_array(18)(315),
      output(19) => mem_array(19)(315),
      output(20) => mem_array(20)(315),
      output(21) => mem_array(21)(315),
      output(22) => mem_array(22)(315),
      output(23) => mem_array(23)(315),
      output(24) => mem_array(24)(315),
      output(25) => mem_array(25)(315),
      output(26) => mem_array(26)(315),
      output(27) => mem_array(27)(315),
      output(28) => mem_array(28)(315),
      output(29) => mem_array(29)(315),
      output(30) => mem_array(30)(315),
      output(31) => mem_array(31)(315),
      output(32) => mem_array(32)(315),
      output(33) => mem_array(33)(315),
      output(34) => mem_array(34)(315),
      output(35) => mem_array(35)(315)
      );
  rom316 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(316),
      output(0)  => mem_array(0)(316),
      output(1)  => mem_array(1)(316),
      output(2)  => mem_array(2)(316),
      output(3)  => mem_array(3)(316),
      output(4)  => mem_array(4)(316),
      output(5)  => mem_array(5)(316),
      output(6)  => mem_array(6)(316),
      output(7)  => mem_array(7)(316),
      output(8)  => mem_array(8)(316),
      output(9)  => mem_array(9)(316),
      output(10) => mem_array(10)(316),
      output(11) => mem_array(11)(316),
      output(12) => mem_array(12)(316),
      output(13) => mem_array(13)(316),
      output(14) => mem_array(14)(316),
      output(15) => mem_array(15)(316),
      output(16) => mem_array(16)(316),
      output(17) => mem_array(17)(316),
      output(18) => mem_array(18)(316),
      output(19) => mem_array(19)(316),
      output(20) => mem_array(20)(316),
      output(21) => mem_array(21)(316),
      output(22) => mem_array(22)(316),
      output(23) => mem_array(23)(316),
      output(24) => mem_array(24)(316),
      output(25) => mem_array(25)(316),
      output(26) => mem_array(26)(316),
      output(27) => mem_array(27)(316),
      output(28) => mem_array(28)(316),
      output(29) => mem_array(29)(316),
      output(30) => mem_array(30)(316),
      output(31) => mem_array(31)(316),
      output(32) => mem_array(32)(316),
      output(33) => mem_array(33)(316),
      output(34) => mem_array(34)(316),
      output(35) => mem_array(35)(316)
      );
  rom317 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(317),
      output(0)  => mem_array(0)(317),
      output(1)  => mem_array(1)(317),
      output(2)  => mem_array(2)(317),
      output(3)  => mem_array(3)(317),
      output(4)  => mem_array(4)(317),
      output(5)  => mem_array(5)(317),
      output(6)  => mem_array(6)(317),
      output(7)  => mem_array(7)(317),
      output(8)  => mem_array(8)(317),
      output(9)  => mem_array(9)(317),
      output(10) => mem_array(10)(317),
      output(11) => mem_array(11)(317),
      output(12) => mem_array(12)(317),
      output(13) => mem_array(13)(317),
      output(14) => mem_array(14)(317),
      output(15) => mem_array(15)(317),
      output(16) => mem_array(16)(317),
      output(17) => mem_array(17)(317),
      output(18) => mem_array(18)(317),
      output(19) => mem_array(19)(317),
      output(20) => mem_array(20)(317),
      output(21) => mem_array(21)(317),
      output(22) => mem_array(22)(317),
      output(23) => mem_array(23)(317),
      output(24) => mem_array(24)(317),
      output(25) => mem_array(25)(317),
      output(26) => mem_array(26)(317),
      output(27) => mem_array(27)(317),
      output(28) => mem_array(28)(317),
      output(29) => mem_array(29)(317),
      output(30) => mem_array(30)(317),
      output(31) => mem_array(31)(317),
      output(32) => mem_array(32)(317),
      output(33) => mem_array(33)(317),
      output(34) => mem_array(34)(317),
      output(35) => mem_array(35)(317)
      );
  rom318 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(318),
      output(0)  => mem_array(0)(318),
      output(1)  => mem_array(1)(318),
      output(2)  => mem_array(2)(318),
      output(3)  => mem_array(3)(318),
      output(4)  => mem_array(4)(318),
      output(5)  => mem_array(5)(318),
      output(6)  => mem_array(6)(318),
      output(7)  => mem_array(7)(318),
      output(8)  => mem_array(8)(318),
      output(9)  => mem_array(9)(318),
      output(10) => mem_array(10)(318),
      output(11) => mem_array(11)(318),
      output(12) => mem_array(12)(318),
      output(13) => mem_array(13)(318),
      output(14) => mem_array(14)(318),
      output(15) => mem_array(15)(318),
      output(16) => mem_array(16)(318),
      output(17) => mem_array(17)(318),
      output(18) => mem_array(18)(318),
      output(19) => mem_array(19)(318),
      output(20) => mem_array(20)(318),
      output(21) => mem_array(21)(318),
      output(22) => mem_array(22)(318),
      output(23) => mem_array(23)(318),
      output(24) => mem_array(24)(318),
      output(25) => mem_array(25)(318),
      output(26) => mem_array(26)(318),
      output(27) => mem_array(27)(318),
      output(28) => mem_array(28)(318),
      output(29) => mem_array(29)(318),
      output(30) => mem_array(30)(318),
      output(31) => mem_array(31)(318),
      output(32) => mem_array(32)(318),
      output(33) => mem_array(33)(318),
      output(34) => mem_array(34)(318),
      output(35) => mem_array(35)(318)
      );
  rom319 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(319),
      output(0)  => mem_array(0)(319),
      output(1)  => mem_array(1)(319),
      output(2)  => mem_array(2)(319),
      output(3)  => mem_array(3)(319),
      output(4)  => mem_array(4)(319),
      output(5)  => mem_array(5)(319),
      output(6)  => mem_array(6)(319),
      output(7)  => mem_array(7)(319),
      output(8)  => mem_array(8)(319),
      output(9)  => mem_array(9)(319),
      output(10) => mem_array(10)(319),
      output(11) => mem_array(11)(319),
      output(12) => mem_array(12)(319),
      output(13) => mem_array(13)(319),
      output(14) => mem_array(14)(319),
      output(15) => mem_array(15)(319),
      output(16) => mem_array(16)(319),
      output(17) => mem_array(17)(319),
      output(18) => mem_array(18)(319),
      output(19) => mem_array(19)(319),
      output(20) => mem_array(20)(319),
      output(21) => mem_array(21)(319),
      output(22) => mem_array(22)(319),
      output(23) => mem_array(23)(319),
      output(24) => mem_array(24)(319),
      output(25) => mem_array(25)(319),
      output(26) => mem_array(26)(319),
      output(27) => mem_array(27)(319),
      output(28) => mem_array(28)(319),
      output(29) => mem_array(29)(319),
      output(30) => mem_array(30)(319),
      output(31) => mem_array(31)(319),
      output(32) => mem_array(32)(319),
      output(33) => mem_array(33)(319),
      output(34) => mem_array(34)(319),
      output(35) => mem_array(35)(319)
      );
  rom320 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(320),
      output(0)  => mem_array(0)(320),
      output(1)  => mem_array(1)(320),
      output(2)  => mem_array(2)(320),
      output(3)  => mem_array(3)(320),
      output(4)  => mem_array(4)(320),
      output(5)  => mem_array(5)(320),
      output(6)  => mem_array(6)(320),
      output(7)  => mem_array(7)(320),
      output(8)  => mem_array(8)(320),
      output(9)  => mem_array(9)(320),
      output(10) => mem_array(10)(320),
      output(11) => mem_array(11)(320),
      output(12) => mem_array(12)(320),
      output(13) => mem_array(13)(320),
      output(14) => mem_array(14)(320),
      output(15) => mem_array(15)(320),
      output(16) => mem_array(16)(320),
      output(17) => mem_array(17)(320),
      output(18) => mem_array(18)(320),
      output(19) => mem_array(19)(320),
      output(20) => mem_array(20)(320),
      output(21) => mem_array(21)(320),
      output(22) => mem_array(22)(320),
      output(23) => mem_array(23)(320),
      output(24) => mem_array(24)(320),
      output(25) => mem_array(25)(320),
      output(26) => mem_array(26)(320),
      output(27) => mem_array(27)(320),
      output(28) => mem_array(28)(320),
      output(29) => mem_array(29)(320),
      output(30) => mem_array(30)(320),
      output(31) => mem_array(31)(320),
      output(32) => mem_array(32)(320),
      output(33) => mem_array(33)(320),
      output(34) => mem_array(34)(320),
      output(35) => mem_array(35)(320)
      );
  rom321 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(321),
      output(0)  => mem_array(0)(321),
      output(1)  => mem_array(1)(321),
      output(2)  => mem_array(2)(321),
      output(3)  => mem_array(3)(321),
      output(4)  => mem_array(4)(321),
      output(5)  => mem_array(5)(321),
      output(6)  => mem_array(6)(321),
      output(7)  => mem_array(7)(321),
      output(8)  => mem_array(8)(321),
      output(9)  => mem_array(9)(321),
      output(10) => mem_array(10)(321),
      output(11) => mem_array(11)(321),
      output(12) => mem_array(12)(321),
      output(13) => mem_array(13)(321),
      output(14) => mem_array(14)(321),
      output(15) => mem_array(15)(321),
      output(16) => mem_array(16)(321),
      output(17) => mem_array(17)(321),
      output(18) => mem_array(18)(321),
      output(19) => mem_array(19)(321),
      output(20) => mem_array(20)(321),
      output(21) => mem_array(21)(321),
      output(22) => mem_array(22)(321),
      output(23) => mem_array(23)(321),
      output(24) => mem_array(24)(321),
      output(25) => mem_array(25)(321),
      output(26) => mem_array(26)(321),
      output(27) => mem_array(27)(321),
      output(28) => mem_array(28)(321),
      output(29) => mem_array(29)(321),
      output(30) => mem_array(30)(321),
      output(31) => mem_array(31)(321),
      output(32) => mem_array(32)(321),
      output(33) => mem_array(33)(321),
      output(34) => mem_array(34)(321),
      output(35) => mem_array(35)(321)
      );
  rom322 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(322),
      output(0)  => mem_array(0)(322),
      output(1)  => mem_array(1)(322),
      output(2)  => mem_array(2)(322),
      output(3)  => mem_array(3)(322),
      output(4)  => mem_array(4)(322),
      output(5)  => mem_array(5)(322),
      output(6)  => mem_array(6)(322),
      output(7)  => mem_array(7)(322),
      output(8)  => mem_array(8)(322),
      output(9)  => mem_array(9)(322),
      output(10) => mem_array(10)(322),
      output(11) => mem_array(11)(322),
      output(12) => mem_array(12)(322),
      output(13) => mem_array(13)(322),
      output(14) => mem_array(14)(322),
      output(15) => mem_array(15)(322),
      output(16) => mem_array(16)(322),
      output(17) => mem_array(17)(322),
      output(18) => mem_array(18)(322),
      output(19) => mem_array(19)(322),
      output(20) => mem_array(20)(322),
      output(21) => mem_array(21)(322),
      output(22) => mem_array(22)(322),
      output(23) => mem_array(23)(322),
      output(24) => mem_array(24)(322),
      output(25) => mem_array(25)(322),
      output(26) => mem_array(26)(322),
      output(27) => mem_array(27)(322),
      output(28) => mem_array(28)(322),
      output(29) => mem_array(29)(322),
      output(30) => mem_array(30)(322),
      output(31) => mem_array(31)(322),
      output(32) => mem_array(32)(322),
      output(33) => mem_array(33)(322),
      output(34) => mem_array(34)(322),
      output(35) => mem_array(35)(322)
      );
  rom323 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(323),
      output(0)  => mem_array(0)(323),
      output(1)  => mem_array(1)(323),
      output(2)  => mem_array(2)(323),
      output(3)  => mem_array(3)(323),
      output(4)  => mem_array(4)(323),
      output(5)  => mem_array(5)(323),
      output(6)  => mem_array(6)(323),
      output(7)  => mem_array(7)(323),
      output(8)  => mem_array(8)(323),
      output(9)  => mem_array(9)(323),
      output(10) => mem_array(10)(323),
      output(11) => mem_array(11)(323),
      output(12) => mem_array(12)(323),
      output(13) => mem_array(13)(323),
      output(14) => mem_array(14)(323),
      output(15) => mem_array(15)(323),
      output(16) => mem_array(16)(323),
      output(17) => mem_array(17)(323),
      output(18) => mem_array(18)(323),
      output(19) => mem_array(19)(323),
      output(20) => mem_array(20)(323),
      output(21) => mem_array(21)(323),
      output(22) => mem_array(22)(323),
      output(23) => mem_array(23)(323),
      output(24) => mem_array(24)(323),
      output(25) => mem_array(25)(323),
      output(26) => mem_array(26)(323),
      output(27) => mem_array(27)(323),
      output(28) => mem_array(28)(323),
      output(29) => mem_array(29)(323),
      output(30) => mem_array(30)(323),
      output(31) => mem_array(31)(323),
      output(32) => mem_array(32)(323),
      output(33) => mem_array(33)(323),
      output(34) => mem_array(34)(323),
      output(35) => mem_array(35)(323)
      );
  rom324 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(324),
      output(0)  => mem_array(0)(324),
      output(1)  => mem_array(1)(324),
      output(2)  => mem_array(2)(324),
      output(3)  => mem_array(3)(324),
      output(4)  => mem_array(4)(324),
      output(5)  => mem_array(5)(324),
      output(6)  => mem_array(6)(324),
      output(7)  => mem_array(7)(324),
      output(8)  => mem_array(8)(324),
      output(9)  => mem_array(9)(324),
      output(10) => mem_array(10)(324),
      output(11) => mem_array(11)(324),
      output(12) => mem_array(12)(324),
      output(13) => mem_array(13)(324),
      output(14) => mem_array(14)(324),
      output(15) => mem_array(15)(324),
      output(16) => mem_array(16)(324),
      output(17) => mem_array(17)(324),
      output(18) => mem_array(18)(324),
      output(19) => mem_array(19)(324),
      output(20) => mem_array(20)(324),
      output(21) => mem_array(21)(324),
      output(22) => mem_array(22)(324),
      output(23) => mem_array(23)(324),
      output(24) => mem_array(24)(324),
      output(25) => mem_array(25)(324),
      output(26) => mem_array(26)(324),
      output(27) => mem_array(27)(324),
      output(28) => mem_array(28)(324),
      output(29) => mem_array(29)(324),
      output(30) => mem_array(30)(324),
      output(31) => mem_array(31)(324),
      output(32) => mem_array(32)(324),
      output(33) => mem_array(33)(324),
      output(34) => mem_array(34)(324),
      output(35) => mem_array(35)(324)
      );
  rom325 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(325),
      output(0)  => mem_array(0)(325),
      output(1)  => mem_array(1)(325),
      output(2)  => mem_array(2)(325),
      output(3)  => mem_array(3)(325),
      output(4)  => mem_array(4)(325),
      output(5)  => mem_array(5)(325),
      output(6)  => mem_array(6)(325),
      output(7)  => mem_array(7)(325),
      output(8)  => mem_array(8)(325),
      output(9)  => mem_array(9)(325),
      output(10) => mem_array(10)(325),
      output(11) => mem_array(11)(325),
      output(12) => mem_array(12)(325),
      output(13) => mem_array(13)(325),
      output(14) => mem_array(14)(325),
      output(15) => mem_array(15)(325),
      output(16) => mem_array(16)(325),
      output(17) => mem_array(17)(325),
      output(18) => mem_array(18)(325),
      output(19) => mem_array(19)(325),
      output(20) => mem_array(20)(325),
      output(21) => mem_array(21)(325),
      output(22) => mem_array(22)(325),
      output(23) => mem_array(23)(325),
      output(24) => mem_array(24)(325),
      output(25) => mem_array(25)(325),
      output(26) => mem_array(26)(325),
      output(27) => mem_array(27)(325),
      output(28) => mem_array(28)(325),
      output(29) => mem_array(29)(325),
      output(30) => mem_array(30)(325),
      output(31) => mem_array(31)(325),
      output(32) => mem_array(32)(325),
      output(33) => mem_array(33)(325),
      output(34) => mem_array(34)(325),
      output(35) => mem_array(35)(325)
      );
  rom326 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(326),
      output(0)  => mem_array(0)(326),
      output(1)  => mem_array(1)(326),
      output(2)  => mem_array(2)(326),
      output(3)  => mem_array(3)(326),
      output(4)  => mem_array(4)(326),
      output(5)  => mem_array(5)(326),
      output(6)  => mem_array(6)(326),
      output(7)  => mem_array(7)(326),
      output(8)  => mem_array(8)(326),
      output(9)  => mem_array(9)(326),
      output(10) => mem_array(10)(326),
      output(11) => mem_array(11)(326),
      output(12) => mem_array(12)(326),
      output(13) => mem_array(13)(326),
      output(14) => mem_array(14)(326),
      output(15) => mem_array(15)(326),
      output(16) => mem_array(16)(326),
      output(17) => mem_array(17)(326),
      output(18) => mem_array(18)(326),
      output(19) => mem_array(19)(326),
      output(20) => mem_array(20)(326),
      output(21) => mem_array(21)(326),
      output(22) => mem_array(22)(326),
      output(23) => mem_array(23)(326),
      output(24) => mem_array(24)(326),
      output(25) => mem_array(25)(326),
      output(26) => mem_array(26)(326),
      output(27) => mem_array(27)(326),
      output(28) => mem_array(28)(326),
      output(29) => mem_array(29)(326),
      output(30) => mem_array(30)(326),
      output(31) => mem_array(31)(326),
      output(32) => mem_array(32)(326),
      output(33) => mem_array(33)(326),
      output(34) => mem_array(34)(326),
      output(35) => mem_array(35)(326)
      );
  rom327 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(327),
      output(0)  => mem_array(0)(327),
      output(1)  => mem_array(1)(327),
      output(2)  => mem_array(2)(327),
      output(3)  => mem_array(3)(327),
      output(4)  => mem_array(4)(327),
      output(5)  => mem_array(5)(327),
      output(6)  => mem_array(6)(327),
      output(7)  => mem_array(7)(327),
      output(8)  => mem_array(8)(327),
      output(9)  => mem_array(9)(327),
      output(10) => mem_array(10)(327),
      output(11) => mem_array(11)(327),
      output(12) => mem_array(12)(327),
      output(13) => mem_array(13)(327),
      output(14) => mem_array(14)(327),
      output(15) => mem_array(15)(327),
      output(16) => mem_array(16)(327),
      output(17) => mem_array(17)(327),
      output(18) => mem_array(18)(327),
      output(19) => mem_array(19)(327),
      output(20) => mem_array(20)(327),
      output(21) => mem_array(21)(327),
      output(22) => mem_array(22)(327),
      output(23) => mem_array(23)(327),
      output(24) => mem_array(24)(327),
      output(25) => mem_array(25)(327),
      output(26) => mem_array(26)(327),
      output(27) => mem_array(27)(327),
      output(28) => mem_array(28)(327),
      output(29) => mem_array(29)(327),
      output(30) => mem_array(30)(327),
      output(31) => mem_array(31)(327),
      output(32) => mem_array(32)(327),
      output(33) => mem_array(33)(327),
      output(34) => mem_array(34)(327),
      output(35) => mem_array(35)(327)
      );
  rom328 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(328),
      output(0)  => mem_array(0)(328),
      output(1)  => mem_array(1)(328),
      output(2)  => mem_array(2)(328),
      output(3)  => mem_array(3)(328),
      output(4)  => mem_array(4)(328),
      output(5)  => mem_array(5)(328),
      output(6)  => mem_array(6)(328),
      output(7)  => mem_array(7)(328),
      output(8)  => mem_array(8)(328),
      output(9)  => mem_array(9)(328),
      output(10) => mem_array(10)(328),
      output(11) => mem_array(11)(328),
      output(12) => mem_array(12)(328),
      output(13) => mem_array(13)(328),
      output(14) => mem_array(14)(328),
      output(15) => mem_array(15)(328),
      output(16) => mem_array(16)(328),
      output(17) => mem_array(17)(328),
      output(18) => mem_array(18)(328),
      output(19) => mem_array(19)(328),
      output(20) => mem_array(20)(328),
      output(21) => mem_array(21)(328),
      output(22) => mem_array(22)(328),
      output(23) => mem_array(23)(328),
      output(24) => mem_array(24)(328),
      output(25) => mem_array(25)(328),
      output(26) => mem_array(26)(328),
      output(27) => mem_array(27)(328),
      output(28) => mem_array(28)(328),
      output(29) => mem_array(29)(328),
      output(30) => mem_array(30)(328),
      output(31) => mem_array(31)(328),
      output(32) => mem_array(32)(328),
      output(33) => mem_array(33)(328),
      output(34) => mem_array(34)(328),
      output(35) => mem_array(35)(328)
      );
  rom329 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(329),
      output(0)  => mem_array(0)(329),
      output(1)  => mem_array(1)(329),
      output(2)  => mem_array(2)(329),
      output(3)  => mem_array(3)(329),
      output(4)  => mem_array(4)(329),
      output(5)  => mem_array(5)(329),
      output(6)  => mem_array(6)(329),
      output(7)  => mem_array(7)(329),
      output(8)  => mem_array(8)(329),
      output(9)  => mem_array(9)(329),
      output(10) => mem_array(10)(329),
      output(11) => mem_array(11)(329),
      output(12) => mem_array(12)(329),
      output(13) => mem_array(13)(329),
      output(14) => mem_array(14)(329),
      output(15) => mem_array(15)(329),
      output(16) => mem_array(16)(329),
      output(17) => mem_array(17)(329),
      output(18) => mem_array(18)(329),
      output(19) => mem_array(19)(329),
      output(20) => mem_array(20)(329),
      output(21) => mem_array(21)(329),
      output(22) => mem_array(22)(329),
      output(23) => mem_array(23)(329),
      output(24) => mem_array(24)(329),
      output(25) => mem_array(25)(329),
      output(26) => mem_array(26)(329),
      output(27) => mem_array(27)(329),
      output(28) => mem_array(28)(329),
      output(29) => mem_array(29)(329),
      output(30) => mem_array(30)(329),
      output(31) => mem_array(31)(329),
      output(32) => mem_array(32)(329),
      output(33) => mem_array(33)(329),
      output(34) => mem_array(34)(329),
      output(35) => mem_array(35)(329)
      );
  rom330 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(330),
      output(0)  => mem_array(0)(330),
      output(1)  => mem_array(1)(330),
      output(2)  => mem_array(2)(330),
      output(3)  => mem_array(3)(330),
      output(4)  => mem_array(4)(330),
      output(5)  => mem_array(5)(330),
      output(6)  => mem_array(6)(330),
      output(7)  => mem_array(7)(330),
      output(8)  => mem_array(8)(330),
      output(9)  => mem_array(9)(330),
      output(10) => mem_array(10)(330),
      output(11) => mem_array(11)(330),
      output(12) => mem_array(12)(330),
      output(13) => mem_array(13)(330),
      output(14) => mem_array(14)(330),
      output(15) => mem_array(15)(330),
      output(16) => mem_array(16)(330),
      output(17) => mem_array(17)(330),
      output(18) => mem_array(18)(330),
      output(19) => mem_array(19)(330),
      output(20) => mem_array(20)(330),
      output(21) => mem_array(21)(330),
      output(22) => mem_array(22)(330),
      output(23) => mem_array(23)(330),
      output(24) => mem_array(24)(330),
      output(25) => mem_array(25)(330),
      output(26) => mem_array(26)(330),
      output(27) => mem_array(27)(330),
      output(28) => mem_array(28)(330),
      output(29) => mem_array(29)(330),
      output(30) => mem_array(30)(330),
      output(31) => mem_array(31)(330),
      output(32) => mem_array(32)(330),
      output(33) => mem_array(33)(330),
      output(34) => mem_array(34)(330),
      output(35) => mem_array(35)(330)
      );
  rom331 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(331),
      output(0)  => mem_array(0)(331),
      output(1)  => mem_array(1)(331),
      output(2)  => mem_array(2)(331),
      output(3)  => mem_array(3)(331),
      output(4)  => mem_array(4)(331),
      output(5)  => mem_array(5)(331),
      output(6)  => mem_array(6)(331),
      output(7)  => mem_array(7)(331),
      output(8)  => mem_array(8)(331),
      output(9)  => mem_array(9)(331),
      output(10) => mem_array(10)(331),
      output(11) => mem_array(11)(331),
      output(12) => mem_array(12)(331),
      output(13) => mem_array(13)(331),
      output(14) => mem_array(14)(331),
      output(15) => mem_array(15)(331),
      output(16) => mem_array(16)(331),
      output(17) => mem_array(17)(331),
      output(18) => mem_array(18)(331),
      output(19) => mem_array(19)(331),
      output(20) => mem_array(20)(331),
      output(21) => mem_array(21)(331),
      output(22) => mem_array(22)(331),
      output(23) => mem_array(23)(331),
      output(24) => mem_array(24)(331),
      output(25) => mem_array(25)(331),
      output(26) => mem_array(26)(331),
      output(27) => mem_array(27)(331),
      output(28) => mem_array(28)(331),
      output(29) => mem_array(29)(331),
      output(30) => mem_array(30)(331),
      output(31) => mem_array(31)(331),
      output(32) => mem_array(32)(331),
      output(33) => mem_array(33)(331),
      output(34) => mem_array(34)(331),
      output(35) => mem_array(35)(331)
      );
  rom332 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(332),
      output(0)  => mem_array(0)(332),
      output(1)  => mem_array(1)(332),
      output(2)  => mem_array(2)(332),
      output(3)  => mem_array(3)(332),
      output(4)  => mem_array(4)(332),
      output(5)  => mem_array(5)(332),
      output(6)  => mem_array(6)(332),
      output(7)  => mem_array(7)(332),
      output(8)  => mem_array(8)(332),
      output(9)  => mem_array(9)(332),
      output(10) => mem_array(10)(332),
      output(11) => mem_array(11)(332),
      output(12) => mem_array(12)(332),
      output(13) => mem_array(13)(332),
      output(14) => mem_array(14)(332),
      output(15) => mem_array(15)(332),
      output(16) => mem_array(16)(332),
      output(17) => mem_array(17)(332),
      output(18) => mem_array(18)(332),
      output(19) => mem_array(19)(332),
      output(20) => mem_array(20)(332),
      output(21) => mem_array(21)(332),
      output(22) => mem_array(22)(332),
      output(23) => mem_array(23)(332),
      output(24) => mem_array(24)(332),
      output(25) => mem_array(25)(332),
      output(26) => mem_array(26)(332),
      output(27) => mem_array(27)(332),
      output(28) => mem_array(28)(332),
      output(29) => mem_array(29)(332),
      output(30) => mem_array(30)(332),
      output(31) => mem_array(31)(332),
      output(32) => mem_array(32)(332),
      output(33) => mem_array(33)(332),
      output(34) => mem_array(34)(332),
      output(35) => mem_array(35)(332)
      );
  rom333 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(333),
      output(0)  => mem_array(0)(333),
      output(1)  => mem_array(1)(333),
      output(2)  => mem_array(2)(333),
      output(3)  => mem_array(3)(333),
      output(4)  => mem_array(4)(333),
      output(5)  => mem_array(5)(333),
      output(6)  => mem_array(6)(333),
      output(7)  => mem_array(7)(333),
      output(8)  => mem_array(8)(333),
      output(9)  => mem_array(9)(333),
      output(10) => mem_array(10)(333),
      output(11) => mem_array(11)(333),
      output(12) => mem_array(12)(333),
      output(13) => mem_array(13)(333),
      output(14) => mem_array(14)(333),
      output(15) => mem_array(15)(333),
      output(16) => mem_array(16)(333),
      output(17) => mem_array(17)(333),
      output(18) => mem_array(18)(333),
      output(19) => mem_array(19)(333),
      output(20) => mem_array(20)(333),
      output(21) => mem_array(21)(333),
      output(22) => mem_array(22)(333),
      output(23) => mem_array(23)(333),
      output(24) => mem_array(24)(333),
      output(25) => mem_array(25)(333),
      output(26) => mem_array(26)(333),
      output(27) => mem_array(27)(333),
      output(28) => mem_array(28)(333),
      output(29) => mem_array(29)(333),
      output(30) => mem_array(30)(333),
      output(31) => mem_array(31)(333),
      output(32) => mem_array(32)(333),
      output(33) => mem_array(33)(333),
      output(34) => mem_array(34)(333),
      output(35) => mem_array(35)(333)
      );
  rom334 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(334),
      output(0)  => mem_array(0)(334),
      output(1)  => mem_array(1)(334),
      output(2)  => mem_array(2)(334),
      output(3)  => mem_array(3)(334),
      output(4)  => mem_array(4)(334),
      output(5)  => mem_array(5)(334),
      output(6)  => mem_array(6)(334),
      output(7)  => mem_array(7)(334),
      output(8)  => mem_array(8)(334),
      output(9)  => mem_array(9)(334),
      output(10) => mem_array(10)(334),
      output(11) => mem_array(11)(334),
      output(12) => mem_array(12)(334),
      output(13) => mem_array(13)(334),
      output(14) => mem_array(14)(334),
      output(15) => mem_array(15)(334),
      output(16) => mem_array(16)(334),
      output(17) => mem_array(17)(334),
      output(18) => mem_array(18)(334),
      output(19) => mem_array(19)(334),
      output(20) => mem_array(20)(334),
      output(21) => mem_array(21)(334),
      output(22) => mem_array(22)(334),
      output(23) => mem_array(23)(334),
      output(24) => mem_array(24)(334),
      output(25) => mem_array(25)(334),
      output(26) => mem_array(26)(334),
      output(27) => mem_array(27)(334),
      output(28) => mem_array(28)(334),
      output(29) => mem_array(29)(334),
      output(30) => mem_array(30)(334),
      output(31) => mem_array(31)(334),
      output(32) => mem_array(32)(334),
      output(33) => mem_array(33)(334),
      output(34) => mem_array(34)(334),
      output(35) => mem_array(35)(334)
      );
  rom335 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(335),
      output(0)  => mem_array(0)(335),
      output(1)  => mem_array(1)(335),
      output(2)  => mem_array(2)(335),
      output(3)  => mem_array(3)(335),
      output(4)  => mem_array(4)(335),
      output(5)  => mem_array(5)(335),
      output(6)  => mem_array(6)(335),
      output(7)  => mem_array(7)(335),
      output(8)  => mem_array(8)(335),
      output(9)  => mem_array(9)(335),
      output(10) => mem_array(10)(335),
      output(11) => mem_array(11)(335),
      output(12) => mem_array(12)(335),
      output(13) => mem_array(13)(335),
      output(14) => mem_array(14)(335),
      output(15) => mem_array(15)(335),
      output(16) => mem_array(16)(335),
      output(17) => mem_array(17)(335),
      output(18) => mem_array(18)(335),
      output(19) => mem_array(19)(335),
      output(20) => mem_array(20)(335),
      output(21) => mem_array(21)(335),
      output(22) => mem_array(22)(335),
      output(23) => mem_array(23)(335),
      output(24) => mem_array(24)(335),
      output(25) => mem_array(25)(335),
      output(26) => mem_array(26)(335),
      output(27) => mem_array(27)(335),
      output(28) => mem_array(28)(335),
      output(29) => mem_array(29)(335),
      output(30) => mem_array(30)(335),
      output(31) => mem_array(31)(335),
      output(32) => mem_array(32)(335),
      output(33) => mem_array(33)(335),
      output(34) => mem_array(34)(335),
      output(35) => mem_array(35)(335)
      );
  rom336 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(336),
      output(0)  => mem_array(0)(336),
      output(1)  => mem_array(1)(336),
      output(2)  => mem_array(2)(336),
      output(3)  => mem_array(3)(336),
      output(4)  => mem_array(4)(336),
      output(5)  => mem_array(5)(336),
      output(6)  => mem_array(6)(336),
      output(7)  => mem_array(7)(336),
      output(8)  => mem_array(8)(336),
      output(9)  => mem_array(9)(336),
      output(10) => mem_array(10)(336),
      output(11) => mem_array(11)(336),
      output(12) => mem_array(12)(336),
      output(13) => mem_array(13)(336),
      output(14) => mem_array(14)(336),
      output(15) => mem_array(15)(336),
      output(16) => mem_array(16)(336),
      output(17) => mem_array(17)(336),
      output(18) => mem_array(18)(336),
      output(19) => mem_array(19)(336),
      output(20) => mem_array(20)(336),
      output(21) => mem_array(21)(336),
      output(22) => mem_array(22)(336),
      output(23) => mem_array(23)(336),
      output(24) => mem_array(24)(336),
      output(25) => mem_array(25)(336),
      output(26) => mem_array(26)(336),
      output(27) => mem_array(27)(336),
      output(28) => mem_array(28)(336),
      output(29) => mem_array(29)(336),
      output(30) => mem_array(30)(336),
      output(31) => mem_array(31)(336),
      output(32) => mem_array(32)(336),
      output(33) => mem_array(33)(336),
      output(34) => mem_array(34)(336),
      output(35) => mem_array(35)(336)
      );
  rom337 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(337),
      output(0)  => mem_array(0)(337),
      output(1)  => mem_array(1)(337),
      output(2)  => mem_array(2)(337),
      output(3)  => mem_array(3)(337),
      output(4)  => mem_array(4)(337),
      output(5)  => mem_array(5)(337),
      output(6)  => mem_array(6)(337),
      output(7)  => mem_array(7)(337),
      output(8)  => mem_array(8)(337),
      output(9)  => mem_array(9)(337),
      output(10) => mem_array(10)(337),
      output(11) => mem_array(11)(337),
      output(12) => mem_array(12)(337),
      output(13) => mem_array(13)(337),
      output(14) => mem_array(14)(337),
      output(15) => mem_array(15)(337),
      output(16) => mem_array(16)(337),
      output(17) => mem_array(17)(337),
      output(18) => mem_array(18)(337),
      output(19) => mem_array(19)(337),
      output(20) => mem_array(20)(337),
      output(21) => mem_array(21)(337),
      output(22) => mem_array(22)(337),
      output(23) => mem_array(23)(337),
      output(24) => mem_array(24)(337),
      output(25) => mem_array(25)(337),
      output(26) => mem_array(26)(337),
      output(27) => mem_array(27)(337),
      output(28) => mem_array(28)(337),
      output(29) => mem_array(29)(337),
      output(30) => mem_array(30)(337),
      output(31) => mem_array(31)(337),
      output(32) => mem_array(32)(337),
      output(33) => mem_array(33)(337),
      output(34) => mem_array(34)(337),
      output(35) => mem_array(35)(337)
      );
  rom338 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(338),
      output(0)  => mem_array(0)(338),
      output(1)  => mem_array(1)(338),
      output(2)  => mem_array(2)(338),
      output(3)  => mem_array(3)(338),
      output(4)  => mem_array(4)(338),
      output(5)  => mem_array(5)(338),
      output(6)  => mem_array(6)(338),
      output(7)  => mem_array(7)(338),
      output(8)  => mem_array(8)(338),
      output(9)  => mem_array(9)(338),
      output(10) => mem_array(10)(338),
      output(11) => mem_array(11)(338),
      output(12) => mem_array(12)(338),
      output(13) => mem_array(13)(338),
      output(14) => mem_array(14)(338),
      output(15) => mem_array(15)(338),
      output(16) => mem_array(16)(338),
      output(17) => mem_array(17)(338),
      output(18) => mem_array(18)(338),
      output(19) => mem_array(19)(338),
      output(20) => mem_array(20)(338),
      output(21) => mem_array(21)(338),
      output(22) => mem_array(22)(338),
      output(23) => mem_array(23)(338),
      output(24) => mem_array(24)(338),
      output(25) => mem_array(25)(338),
      output(26) => mem_array(26)(338),
      output(27) => mem_array(27)(338),
      output(28) => mem_array(28)(338),
      output(29) => mem_array(29)(338),
      output(30) => mem_array(30)(338),
      output(31) => mem_array(31)(338),
      output(32) => mem_array(32)(338),
      output(33) => mem_array(33)(338),
      output(34) => mem_array(34)(338),
      output(35) => mem_array(35)(338)
      );
  rom339 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(339),
      output(0)  => mem_array(0)(339),
      output(1)  => mem_array(1)(339),
      output(2)  => mem_array(2)(339),
      output(3)  => mem_array(3)(339),
      output(4)  => mem_array(4)(339),
      output(5)  => mem_array(5)(339),
      output(6)  => mem_array(6)(339),
      output(7)  => mem_array(7)(339),
      output(8)  => mem_array(8)(339),
      output(9)  => mem_array(9)(339),
      output(10) => mem_array(10)(339),
      output(11) => mem_array(11)(339),
      output(12) => mem_array(12)(339),
      output(13) => mem_array(13)(339),
      output(14) => mem_array(14)(339),
      output(15) => mem_array(15)(339),
      output(16) => mem_array(16)(339),
      output(17) => mem_array(17)(339),
      output(18) => mem_array(18)(339),
      output(19) => mem_array(19)(339),
      output(20) => mem_array(20)(339),
      output(21) => mem_array(21)(339),
      output(22) => mem_array(22)(339),
      output(23) => mem_array(23)(339),
      output(24) => mem_array(24)(339),
      output(25) => mem_array(25)(339),
      output(26) => mem_array(26)(339),
      output(27) => mem_array(27)(339),
      output(28) => mem_array(28)(339),
      output(29) => mem_array(29)(339),
      output(30) => mem_array(30)(339),
      output(31) => mem_array(31)(339),
      output(32) => mem_array(32)(339),
      output(33) => mem_array(33)(339),
      output(34) => mem_array(34)(339),
      output(35) => mem_array(35)(339)
      );
  rom340 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(340),
      output(0)  => mem_array(0)(340),
      output(1)  => mem_array(1)(340),
      output(2)  => mem_array(2)(340),
      output(3)  => mem_array(3)(340),
      output(4)  => mem_array(4)(340),
      output(5)  => mem_array(5)(340),
      output(6)  => mem_array(6)(340),
      output(7)  => mem_array(7)(340),
      output(8)  => mem_array(8)(340),
      output(9)  => mem_array(9)(340),
      output(10) => mem_array(10)(340),
      output(11) => mem_array(11)(340),
      output(12) => mem_array(12)(340),
      output(13) => mem_array(13)(340),
      output(14) => mem_array(14)(340),
      output(15) => mem_array(15)(340),
      output(16) => mem_array(16)(340),
      output(17) => mem_array(17)(340),
      output(18) => mem_array(18)(340),
      output(19) => mem_array(19)(340),
      output(20) => mem_array(20)(340),
      output(21) => mem_array(21)(340),
      output(22) => mem_array(22)(340),
      output(23) => mem_array(23)(340),
      output(24) => mem_array(24)(340),
      output(25) => mem_array(25)(340),
      output(26) => mem_array(26)(340),
      output(27) => mem_array(27)(340),
      output(28) => mem_array(28)(340),
      output(29) => mem_array(29)(340),
      output(30) => mem_array(30)(340),
      output(31) => mem_array(31)(340),
      output(32) => mem_array(32)(340),
      output(33) => mem_array(33)(340),
      output(34) => mem_array(34)(340),
      output(35) => mem_array(35)(340)
      );
  rom341 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(341),
      output(0)  => mem_array(0)(341),
      output(1)  => mem_array(1)(341),
      output(2)  => mem_array(2)(341),
      output(3)  => mem_array(3)(341),
      output(4)  => mem_array(4)(341),
      output(5)  => mem_array(5)(341),
      output(6)  => mem_array(6)(341),
      output(7)  => mem_array(7)(341),
      output(8)  => mem_array(8)(341),
      output(9)  => mem_array(9)(341),
      output(10) => mem_array(10)(341),
      output(11) => mem_array(11)(341),
      output(12) => mem_array(12)(341),
      output(13) => mem_array(13)(341),
      output(14) => mem_array(14)(341),
      output(15) => mem_array(15)(341),
      output(16) => mem_array(16)(341),
      output(17) => mem_array(17)(341),
      output(18) => mem_array(18)(341),
      output(19) => mem_array(19)(341),
      output(20) => mem_array(20)(341),
      output(21) => mem_array(21)(341),
      output(22) => mem_array(22)(341),
      output(23) => mem_array(23)(341),
      output(24) => mem_array(24)(341),
      output(25) => mem_array(25)(341),
      output(26) => mem_array(26)(341),
      output(27) => mem_array(27)(341),
      output(28) => mem_array(28)(341),
      output(29) => mem_array(29)(341),
      output(30) => mem_array(30)(341),
      output(31) => mem_array(31)(341),
      output(32) => mem_array(32)(341),
      output(33) => mem_array(33)(341),
      output(34) => mem_array(34)(341),
      output(35) => mem_array(35)(341)
      );
  rom342 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(342),
      output(0)  => mem_array(0)(342),
      output(1)  => mem_array(1)(342),
      output(2)  => mem_array(2)(342),
      output(3)  => mem_array(3)(342),
      output(4)  => mem_array(4)(342),
      output(5)  => mem_array(5)(342),
      output(6)  => mem_array(6)(342),
      output(7)  => mem_array(7)(342),
      output(8)  => mem_array(8)(342),
      output(9)  => mem_array(9)(342),
      output(10) => mem_array(10)(342),
      output(11) => mem_array(11)(342),
      output(12) => mem_array(12)(342),
      output(13) => mem_array(13)(342),
      output(14) => mem_array(14)(342),
      output(15) => mem_array(15)(342),
      output(16) => mem_array(16)(342),
      output(17) => mem_array(17)(342),
      output(18) => mem_array(18)(342),
      output(19) => mem_array(19)(342),
      output(20) => mem_array(20)(342),
      output(21) => mem_array(21)(342),
      output(22) => mem_array(22)(342),
      output(23) => mem_array(23)(342),
      output(24) => mem_array(24)(342),
      output(25) => mem_array(25)(342),
      output(26) => mem_array(26)(342),
      output(27) => mem_array(27)(342),
      output(28) => mem_array(28)(342),
      output(29) => mem_array(29)(342),
      output(30) => mem_array(30)(342),
      output(31) => mem_array(31)(342),
      output(32) => mem_array(32)(342),
      output(33) => mem_array(33)(342),
      output(34) => mem_array(34)(342),
      output(35) => mem_array(35)(342)
      );
  rom343 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(343),
      output(0)  => mem_array(0)(343),
      output(1)  => mem_array(1)(343),
      output(2)  => mem_array(2)(343),
      output(3)  => mem_array(3)(343),
      output(4)  => mem_array(4)(343),
      output(5)  => mem_array(5)(343),
      output(6)  => mem_array(6)(343),
      output(7)  => mem_array(7)(343),
      output(8)  => mem_array(8)(343),
      output(9)  => mem_array(9)(343),
      output(10) => mem_array(10)(343),
      output(11) => mem_array(11)(343),
      output(12) => mem_array(12)(343),
      output(13) => mem_array(13)(343),
      output(14) => mem_array(14)(343),
      output(15) => mem_array(15)(343),
      output(16) => mem_array(16)(343),
      output(17) => mem_array(17)(343),
      output(18) => mem_array(18)(343),
      output(19) => mem_array(19)(343),
      output(20) => mem_array(20)(343),
      output(21) => mem_array(21)(343),
      output(22) => mem_array(22)(343),
      output(23) => mem_array(23)(343),
      output(24) => mem_array(24)(343),
      output(25) => mem_array(25)(343),
      output(26) => mem_array(26)(343),
      output(27) => mem_array(27)(343),
      output(28) => mem_array(28)(343),
      output(29) => mem_array(29)(343),
      output(30) => mem_array(30)(343),
      output(31) => mem_array(31)(343),
      output(32) => mem_array(32)(343),
      output(33) => mem_array(33)(343),
      output(34) => mem_array(34)(343),
      output(35) => mem_array(35)(343)
      );
  rom344 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(344),
      output(0)  => mem_array(0)(344),
      output(1)  => mem_array(1)(344),
      output(2)  => mem_array(2)(344),
      output(3)  => mem_array(3)(344),
      output(4)  => mem_array(4)(344),
      output(5)  => mem_array(5)(344),
      output(6)  => mem_array(6)(344),
      output(7)  => mem_array(7)(344),
      output(8)  => mem_array(8)(344),
      output(9)  => mem_array(9)(344),
      output(10) => mem_array(10)(344),
      output(11) => mem_array(11)(344),
      output(12) => mem_array(12)(344),
      output(13) => mem_array(13)(344),
      output(14) => mem_array(14)(344),
      output(15) => mem_array(15)(344),
      output(16) => mem_array(16)(344),
      output(17) => mem_array(17)(344),
      output(18) => mem_array(18)(344),
      output(19) => mem_array(19)(344),
      output(20) => mem_array(20)(344),
      output(21) => mem_array(21)(344),
      output(22) => mem_array(22)(344),
      output(23) => mem_array(23)(344),
      output(24) => mem_array(24)(344),
      output(25) => mem_array(25)(344),
      output(26) => mem_array(26)(344),
      output(27) => mem_array(27)(344),
      output(28) => mem_array(28)(344),
      output(29) => mem_array(29)(344),
      output(30) => mem_array(30)(344),
      output(31) => mem_array(31)(344),
      output(32) => mem_array(32)(344),
      output(33) => mem_array(33)(344),
      output(34) => mem_array(34)(344),
      output(35) => mem_array(35)(344)
      );
  rom345 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000100100000001101010000")
    port map (
      enable_o   => mem_enable_lines(345),
      output(0)  => mem_array(0)(345),
      output(1)  => mem_array(1)(345),
      output(2)  => mem_array(2)(345),
      output(3)  => mem_array(3)(345),
      output(4)  => mem_array(4)(345),
      output(5)  => mem_array(5)(345),
      output(6)  => mem_array(6)(345),
      output(7)  => mem_array(7)(345),
      output(8)  => mem_array(8)(345),
      output(9)  => mem_array(9)(345),
      output(10) => mem_array(10)(345),
      output(11) => mem_array(11)(345),
      output(12) => mem_array(12)(345),
      output(13) => mem_array(13)(345),
      output(14) => mem_array(14)(345),
      output(15) => mem_array(15)(345),
      output(16) => mem_array(16)(345),
      output(17) => mem_array(17)(345),
      output(18) => mem_array(18)(345),
      output(19) => mem_array(19)(345),
      output(20) => mem_array(20)(345),
      output(21) => mem_array(21)(345),
      output(22) => mem_array(22)(345),
      output(23) => mem_array(23)(345),
      output(24) => mem_array(24)(345),
      output(25) => mem_array(25)(345),
      output(26) => mem_array(26)(345),
      output(27) => mem_array(27)(345),
      output(28) => mem_array(28)(345),
      output(29) => mem_array(29)(345),
      output(30) => mem_array(30)(345),
      output(31) => mem_array(31)(345),
      output(32) => mem_array(32)(345),
      output(33) => mem_array(33)(345),
      output(34) => mem_array(34)(345),
      output(35) => mem_array(35)(345)
      );
  rom346 : entity work.rom
    generic map (
      bits  => 36,
      value => "001000010001000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(346),
      output(0)  => mem_array(0)(346),
      output(1)  => mem_array(1)(346),
      output(2)  => mem_array(2)(346),
      output(3)  => mem_array(3)(346),
      output(4)  => mem_array(4)(346),
      output(5)  => mem_array(5)(346),
      output(6)  => mem_array(6)(346),
      output(7)  => mem_array(7)(346),
      output(8)  => mem_array(8)(346),
      output(9)  => mem_array(9)(346),
      output(10) => mem_array(10)(346),
      output(11) => mem_array(11)(346),
      output(12) => mem_array(12)(346),
      output(13) => mem_array(13)(346),
      output(14) => mem_array(14)(346),
      output(15) => mem_array(15)(346),
      output(16) => mem_array(16)(346),
      output(17) => mem_array(17)(346),
      output(18) => mem_array(18)(346),
      output(19) => mem_array(19)(346),
      output(20) => mem_array(20)(346),
      output(21) => mem_array(21)(346),
      output(22) => mem_array(22)(346),
      output(23) => mem_array(23)(346),
      output(24) => mem_array(24)(346),
      output(25) => mem_array(25)(346),
      output(26) => mem_array(26)(346),
      output(27) => mem_array(27)(346),
      output(28) => mem_array(28)(346),
      output(29) => mem_array(29)(346),
      output(30) => mem_array(30)(346),
      output(31) => mem_array(31)(346),
      output(32) => mem_array(32)(346),
      output(33) => mem_array(33)(346),
      output(34) => mem_array(34)(346),
      output(35) => mem_array(35)(346)
      );
  rom347 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(347),
      output(0)  => mem_array(0)(347),
      output(1)  => mem_array(1)(347),
      output(2)  => mem_array(2)(347),
      output(3)  => mem_array(3)(347),
      output(4)  => mem_array(4)(347),
      output(5)  => mem_array(5)(347),
      output(6)  => mem_array(6)(347),
      output(7)  => mem_array(7)(347),
      output(8)  => mem_array(8)(347),
      output(9)  => mem_array(9)(347),
      output(10) => mem_array(10)(347),
      output(11) => mem_array(11)(347),
      output(12) => mem_array(12)(347),
      output(13) => mem_array(13)(347),
      output(14) => mem_array(14)(347),
      output(15) => mem_array(15)(347),
      output(16) => mem_array(16)(347),
      output(17) => mem_array(17)(347),
      output(18) => mem_array(18)(347),
      output(19) => mem_array(19)(347),
      output(20) => mem_array(20)(347),
      output(21) => mem_array(21)(347),
      output(22) => mem_array(22)(347),
      output(23) => mem_array(23)(347),
      output(24) => mem_array(24)(347),
      output(25) => mem_array(25)(347),
      output(26) => mem_array(26)(347),
      output(27) => mem_array(27)(347),
      output(28) => mem_array(28)(347),
      output(29) => mem_array(29)(347),
      output(30) => mem_array(30)(347),
      output(31) => mem_array(31)(347),
      output(32) => mem_array(32)(347),
      output(33) => mem_array(33)(347),
      output(34) => mem_array(34)(347),
      output(35) => mem_array(35)(347)
      );
  rom348 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(348),
      output(0)  => mem_array(0)(348),
      output(1)  => mem_array(1)(348),
      output(2)  => mem_array(2)(348),
      output(3)  => mem_array(3)(348),
      output(4)  => mem_array(4)(348),
      output(5)  => mem_array(5)(348),
      output(6)  => mem_array(6)(348),
      output(7)  => mem_array(7)(348),
      output(8)  => mem_array(8)(348),
      output(9)  => mem_array(9)(348),
      output(10) => mem_array(10)(348),
      output(11) => mem_array(11)(348),
      output(12) => mem_array(12)(348),
      output(13) => mem_array(13)(348),
      output(14) => mem_array(14)(348),
      output(15) => mem_array(15)(348),
      output(16) => mem_array(16)(348),
      output(17) => mem_array(17)(348),
      output(18) => mem_array(18)(348),
      output(19) => mem_array(19)(348),
      output(20) => mem_array(20)(348),
      output(21) => mem_array(21)(348),
      output(22) => mem_array(22)(348),
      output(23) => mem_array(23)(348),
      output(24) => mem_array(24)(348),
      output(25) => mem_array(25)(348),
      output(26) => mem_array(26)(348),
      output(27) => mem_array(27)(348),
      output(28) => mem_array(28)(348),
      output(29) => mem_array(29)(348),
      output(30) => mem_array(30)(348),
      output(31) => mem_array(31)(348),
      output(32) => mem_array(32)(348),
      output(33) => mem_array(33)(348),
      output(34) => mem_array(34)(348),
      output(35) => mem_array(35)(348)
      );
  rom349 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(349),
      output(0)  => mem_array(0)(349),
      output(1)  => mem_array(1)(349),
      output(2)  => mem_array(2)(349),
      output(3)  => mem_array(3)(349),
      output(4)  => mem_array(4)(349),
      output(5)  => mem_array(5)(349),
      output(6)  => mem_array(6)(349),
      output(7)  => mem_array(7)(349),
      output(8)  => mem_array(8)(349),
      output(9)  => mem_array(9)(349),
      output(10) => mem_array(10)(349),
      output(11) => mem_array(11)(349),
      output(12) => mem_array(12)(349),
      output(13) => mem_array(13)(349),
      output(14) => mem_array(14)(349),
      output(15) => mem_array(15)(349),
      output(16) => mem_array(16)(349),
      output(17) => mem_array(17)(349),
      output(18) => mem_array(18)(349),
      output(19) => mem_array(19)(349),
      output(20) => mem_array(20)(349),
      output(21) => mem_array(21)(349),
      output(22) => mem_array(22)(349),
      output(23) => mem_array(23)(349),
      output(24) => mem_array(24)(349),
      output(25) => mem_array(25)(349),
      output(26) => mem_array(26)(349),
      output(27) => mem_array(27)(349),
      output(28) => mem_array(28)(349),
      output(29) => mem_array(29)(349),
      output(30) => mem_array(30)(349),
      output(31) => mem_array(31)(349),
      output(32) => mem_array(32)(349),
      output(33) => mem_array(33)(349),
      output(34) => mem_array(34)(349),
      output(35) => mem_array(35)(349)
      );
  rom350 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(350),
      output(0)  => mem_array(0)(350),
      output(1)  => mem_array(1)(350),
      output(2)  => mem_array(2)(350),
      output(3)  => mem_array(3)(350),
      output(4)  => mem_array(4)(350),
      output(5)  => mem_array(5)(350),
      output(6)  => mem_array(6)(350),
      output(7)  => mem_array(7)(350),
      output(8)  => mem_array(8)(350),
      output(9)  => mem_array(9)(350),
      output(10) => mem_array(10)(350),
      output(11) => mem_array(11)(350),
      output(12) => mem_array(12)(350),
      output(13) => mem_array(13)(350),
      output(14) => mem_array(14)(350),
      output(15) => mem_array(15)(350),
      output(16) => mem_array(16)(350),
      output(17) => mem_array(17)(350),
      output(18) => mem_array(18)(350),
      output(19) => mem_array(19)(350),
      output(20) => mem_array(20)(350),
      output(21) => mem_array(21)(350),
      output(22) => mem_array(22)(350),
      output(23) => mem_array(23)(350),
      output(24) => mem_array(24)(350),
      output(25) => mem_array(25)(350),
      output(26) => mem_array(26)(350),
      output(27) => mem_array(27)(350),
      output(28) => mem_array(28)(350),
      output(29) => mem_array(29)(350),
      output(30) => mem_array(30)(350),
      output(31) => mem_array(31)(350),
      output(32) => mem_array(32)(350),
      output(33) => mem_array(33)(350),
      output(34) => mem_array(34)(350),
      output(35) => mem_array(35)(350)
      );
  rom351 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(351),
      output(0)  => mem_array(0)(351),
      output(1)  => mem_array(1)(351),
      output(2)  => mem_array(2)(351),
      output(3)  => mem_array(3)(351),
      output(4)  => mem_array(4)(351),
      output(5)  => mem_array(5)(351),
      output(6)  => mem_array(6)(351),
      output(7)  => mem_array(7)(351),
      output(8)  => mem_array(8)(351),
      output(9)  => mem_array(9)(351),
      output(10) => mem_array(10)(351),
      output(11) => mem_array(11)(351),
      output(12) => mem_array(12)(351),
      output(13) => mem_array(13)(351),
      output(14) => mem_array(14)(351),
      output(15) => mem_array(15)(351),
      output(16) => mem_array(16)(351),
      output(17) => mem_array(17)(351),
      output(18) => mem_array(18)(351),
      output(19) => mem_array(19)(351),
      output(20) => mem_array(20)(351),
      output(21) => mem_array(21)(351),
      output(22) => mem_array(22)(351),
      output(23) => mem_array(23)(351),
      output(24) => mem_array(24)(351),
      output(25) => mem_array(25)(351),
      output(26) => mem_array(26)(351),
      output(27) => mem_array(27)(351),
      output(28) => mem_array(28)(351),
      output(29) => mem_array(29)(351),
      output(30) => mem_array(30)(351),
      output(31) => mem_array(31)(351),
      output(32) => mem_array(32)(351),
      output(33) => mem_array(33)(351),
      output(34) => mem_array(34)(351),
      output(35) => mem_array(35)(351)
      );
  rom352 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(352),
      output(0)  => mem_array(0)(352),
      output(1)  => mem_array(1)(352),
      output(2)  => mem_array(2)(352),
      output(3)  => mem_array(3)(352),
      output(4)  => mem_array(4)(352),
      output(5)  => mem_array(5)(352),
      output(6)  => mem_array(6)(352),
      output(7)  => mem_array(7)(352),
      output(8)  => mem_array(8)(352),
      output(9)  => mem_array(9)(352),
      output(10) => mem_array(10)(352),
      output(11) => mem_array(11)(352),
      output(12) => mem_array(12)(352),
      output(13) => mem_array(13)(352),
      output(14) => mem_array(14)(352),
      output(15) => mem_array(15)(352),
      output(16) => mem_array(16)(352),
      output(17) => mem_array(17)(352),
      output(18) => mem_array(18)(352),
      output(19) => mem_array(19)(352),
      output(20) => mem_array(20)(352),
      output(21) => mem_array(21)(352),
      output(22) => mem_array(22)(352),
      output(23) => mem_array(23)(352),
      output(24) => mem_array(24)(352),
      output(25) => mem_array(25)(352),
      output(26) => mem_array(26)(352),
      output(27) => mem_array(27)(352),
      output(28) => mem_array(28)(352),
      output(29) => mem_array(29)(352),
      output(30) => mem_array(30)(352),
      output(31) => mem_array(31)(352),
      output(32) => mem_array(32)(352),
      output(33) => mem_array(33)(352),
      output(34) => mem_array(34)(352),
      output(35) => mem_array(35)(352)
      );
  rom353 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(353),
      output(0)  => mem_array(0)(353),
      output(1)  => mem_array(1)(353),
      output(2)  => mem_array(2)(353),
      output(3)  => mem_array(3)(353),
      output(4)  => mem_array(4)(353),
      output(5)  => mem_array(5)(353),
      output(6)  => mem_array(6)(353),
      output(7)  => mem_array(7)(353),
      output(8)  => mem_array(8)(353),
      output(9)  => mem_array(9)(353),
      output(10) => mem_array(10)(353),
      output(11) => mem_array(11)(353),
      output(12) => mem_array(12)(353),
      output(13) => mem_array(13)(353),
      output(14) => mem_array(14)(353),
      output(15) => mem_array(15)(353),
      output(16) => mem_array(16)(353),
      output(17) => mem_array(17)(353),
      output(18) => mem_array(18)(353),
      output(19) => mem_array(19)(353),
      output(20) => mem_array(20)(353),
      output(21) => mem_array(21)(353),
      output(22) => mem_array(22)(353),
      output(23) => mem_array(23)(353),
      output(24) => mem_array(24)(353),
      output(25) => mem_array(25)(353),
      output(26) => mem_array(26)(353),
      output(27) => mem_array(27)(353),
      output(28) => mem_array(28)(353),
      output(29) => mem_array(29)(353),
      output(30) => mem_array(30)(353),
      output(31) => mem_array(31)(353),
      output(32) => mem_array(32)(353),
      output(33) => mem_array(33)(353),
      output(34) => mem_array(34)(353),
      output(35) => mem_array(35)(353)
      );
  rom354 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(354),
      output(0)  => mem_array(0)(354),
      output(1)  => mem_array(1)(354),
      output(2)  => mem_array(2)(354),
      output(3)  => mem_array(3)(354),
      output(4)  => mem_array(4)(354),
      output(5)  => mem_array(5)(354),
      output(6)  => mem_array(6)(354),
      output(7)  => mem_array(7)(354),
      output(8)  => mem_array(8)(354),
      output(9)  => mem_array(9)(354),
      output(10) => mem_array(10)(354),
      output(11) => mem_array(11)(354),
      output(12) => mem_array(12)(354),
      output(13) => mem_array(13)(354),
      output(14) => mem_array(14)(354),
      output(15) => mem_array(15)(354),
      output(16) => mem_array(16)(354),
      output(17) => mem_array(17)(354),
      output(18) => mem_array(18)(354),
      output(19) => mem_array(19)(354),
      output(20) => mem_array(20)(354),
      output(21) => mem_array(21)(354),
      output(22) => mem_array(22)(354),
      output(23) => mem_array(23)(354),
      output(24) => mem_array(24)(354),
      output(25) => mem_array(25)(354),
      output(26) => mem_array(26)(354),
      output(27) => mem_array(27)(354),
      output(28) => mem_array(28)(354),
      output(29) => mem_array(29)(354),
      output(30) => mem_array(30)(354),
      output(31) => mem_array(31)(354),
      output(32) => mem_array(32)(354),
      output(33) => mem_array(33)(354),
      output(34) => mem_array(34)(354),
      output(35) => mem_array(35)(354)
      );
  rom355 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(355),
      output(0)  => mem_array(0)(355),
      output(1)  => mem_array(1)(355),
      output(2)  => mem_array(2)(355),
      output(3)  => mem_array(3)(355),
      output(4)  => mem_array(4)(355),
      output(5)  => mem_array(5)(355),
      output(6)  => mem_array(6)(355),
      output(7)  => mem_array(7)(355),
      output(8)  => mem_array(8)(355),
      output(9)  => mem_array(9)(355),
      output(10) => mem_array(10)(355),
      output(11) => mem_array(11)(355),
      output(12) => mem_array(12)(355),
      output(13) => mem_array(13)(355),
      output(14) => mem_array(14)(355),
      output(15) => mem_array(15)(355),
      output(16) => mem_array(16)(355),
      output(17) => mem_array(17)(355),
      output(18) => mem_array(18)(355),
      output(19) => mem_array(19)(355),
      output(20) => mem_array(20)(355),
      output(21) => mem_array(21)(355),
      output(22) => mem_array(22)(355),
      output(23) => mem_array(23)(355),
      output(24) => mem_array(24)(355),
      output(25) => mem_array(25)(355),
      output(26) => mem_array(26)(355),
      output(27) => mem_array(27)(355),
      output(28) => mem_array(28)(355),
      output(29) => mem_array(29)(355),
      output(30) => mem_array(30)(355),
      output(31) => mem_array(31)(355),
      output(32) => mem_array(32)(355),
      output(33) => mem_array(33)(355),
      output(34) => mem_array(34)(355),
      output(35) => mem_array(35)(355)
      );
  rom356 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(356),
      output(0)  => mem_array(0)(356),
      output(1)  => mem_array(1)(356),
      output(2)  => mem_array(2)(356),
      output(3)  => mem_array(3)(356),
      output(4)  => mem_array(4)(356),
      output(5)  => mem_array(5)(356),
      output(6)  => mem_array(6)(356),
      output(7)  => mem_array(7)(356),
      output(8)  => mem_array(8)(356),
      output(9)  => mem_array(9)(356),
      output(10) => mem_array(10)(356),
      output(11) => mem_array(11)(356),
      output(12) => mem_array(12)(356),
      output(13) => mem_array(13)(356),
      output(14) => mem_array(14)(356),
      output(15) => mem_array(15)(356),
      output(16) => mem_array(16)(356),
      output(17) => mem_array(17)(356),
      output(18) => mem_array(18)(356),
      output(19) => mem_array(19)(356),
      output(20) => mem_array(20)(356),
      output(21) => mem_array(21)(356),
      output(22) => mem_array(22)(356),
      output(23) => mem_array(23)(356),
      output(24) => mem_array(24)(356),
      output(25) => mem_array(25)(356),
      output(26) => mem_array(26)(356),
      output(27) => mem_array(27)(356),
      output(28) => mem_array(28)(356),
      output(29) => mem_array(29)(356),
      output(30) => mem_array(30)(356),
      output(31) => mem_array(31)(356),
      output(32) => mem_array(32)(356),
      output(33) => mem_array(33)(356),
      output(34) => mem_array(34)(356),
      output(35) => mem_array(35)(356)
      );
  rom357 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(357),
      output(0)  => mem_array(0)(357),
      output(1)  => mem_array(1)(357),
      output(2)  => mem_array(2)(357),
      output(3)  => mem_array(3)(357),
      output(4)  => mem_array(4)(357),
      output(5)  => mem_array(5)(357),
      output(6)  => mem_array(6)(357),
      output(7)  => mem_array(7)(357),
      output(8)  => mem_array(8)(357),
      output(9)  => mem_array(9)(357),
      output(10) => mem_array(10)(357),
      output(11) => mem_array(11)(357),
      output(12) => mem_array(12)(357),
      output(13) => mem_array(13)(357),
      output(14) => mem_array(14)(357),
      output(15) => mem_array(15)(357),
      output(16) => mem_array(16)(357),
      output(17) => mem_array(17)(357),
      output(18) => mem_array(18)(357),
      output(19) => mem_array(19)(357),
      output(20) => mem_array(20)(357),
      output(21) => mem_array(21)(357),
      output(22) => mem_array(22)(357),
      output(23) => mem_array(23)(357),
      output(24) => mem_array(24)(357),
      output(25) => mem_array(25)(357),
      output(26) => mem_array(26)(357),
      output(27) => mem_array(27)(357),
      output(28) => mem_array(28)(357),
      output(29) => mem_array(29)(357),
      output(30) => mem_array(30)(357),
      output(31) => mem_array(31)(357),
      output(32) => mem_array(32)(357),
      output(33) => mem_array(33)(357),
      output(34) => mem_array(34)(357),
      output(35) => mem_array(35)(357)
      );
  rom358 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(358),
      output(0)  => mem_array(0)(358),
      output(1)  => mem_array(1)(358),
      output(2)  => mem_array(2)(358),
      output(3)  => mem_array(3)(358),
      output(4)  => mem_array(4)(358),
      output(5)  => mem_array(5)(358),
      output(6)  => mem_array(6)(358),
      output(7)  => mem_array(7)(358),
      output(8)  => mem_array(8)(358),
      output(9)  => mem_array(9)(358),
      output(10) => mem_array(10)(358),
      output(11) => mem_array(11)(358),
      output(12) => mem_array(12)(358),
      output(13) => mem_array(13)(358),
      output(14) => mem_array(14)(358),
      output(15) => mem_array(15)(358),
      output(16) => mem_array(16)(358),
      output(17) => mem_array(17)(358),
      output(18) => mem_array(18)(358),
      output(19) => mem_array(19)(358),
      output(20) => mem_array(20)(358),
      output(21) => mem_array(21)(358),
      output(22) => mem_array(22)(358),
      output(23) => mem_array(23)(358),
      output(24) => mem_array(24)(358),
      output(25) => mem_array(25)(358),
      output(26) => mem_array(26)(358),
      output(27) => mem_array(27)(358),
      output(28) => mem_array(28)(358),
      output(29) => mem_array(29)(358),
      output(30) => mem_array(30)(358),
      output(31) => mem_array(31)(358),
      output(32) => mem_array(32)(358),
      output(33) => mem_array(33)(358),
      output(34) => mem_array(34)(358),
      output(35) => mem_array(35)(358)
      );
  rom359 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(359),
      output(0)  => mem_array(0)(359),
      output(1)  => mem_array(1)(359),
      output(2)  => mem_array(2)(359),
      output(3)  => mem_array(3)(359),
      output(4)  => mem_array(4)(359),
      output(5)  => mem_array(5)(359),
      output(6)  => mem_array(6)(359),
      output(7)  => mem_array(7)(359),
      output(8)  => mem_array(8)(359),
      output(9)  => mem_array(9)(359),
      output(10) => mem_array(10)(359),
      output(11) => mem_array(11)(359),
      output(12) => mem_array(12)(359),
      output(13) => mem_array(13)(359),
      output(14) => mem_array(14)(359),
      output(15) => mem_array(15)(359),
      output(16) => mem_array(16)(359),
      output(17) => mem_array(17)(359),
      output(18) => mem_array(18)(359),
      output(19) => mem_array(19)(359),
      output(20) => mem_array(20)(359),
      output(21) => mem_array(21)(359),
      output(22) => mem_array(22)(359),
      output(23) => mem_array(23)(359),
      output(24) => mem_array(24)(359),
      output(25) => mem_array(25)(359),
      output(26) => mem_array(26)(359),
      output(27) => mem_array(27)(359),
      output(28) => mem_array(28)(359),
      output(29) => mem_array(29)(359),
      output(30) => mem_array(30)(359),
      output(31) => mem_array(31)(359),
      output(32) => mem_array(32)(359),
      output(33) => mem_array(33)(359),
      output(34) => mem_array(34)(359),
      output(35) => mem_array(35)(359)
      );
  rom360 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(360),
      output(0)  => mem_array(0)(360),
      output(1)  => mem_array(1)(360),
      output(2)  => mem_array(2)(360),
      output(3)  => mem_array(3)(360),
      output(4)  => mem_array(4)(360),
      output(5)  => mem_array(5)(360),
      output(6)  => mem_array(6)(360),
      output(7)  => mem_array(7)(360),
      output(8)  => mem_array(8)(360),
      output(9)  => mem_array(9)(360),
      output(10) => mem_array(10)(360),
      output(11) => mem_array(11)(360),
      output(12) => mem_array(12)(360),
      output(13) => mem_array(13)(360),
      output(14) => mem_array(14)(360),
      output(15) => mem_array(15)(360),
      output(16) => mem_array(16)(360),
      output(17) => mem_array(17)(360),
      output(18) => mem_array(18)(360),
      output(19) => mem_array(19)(360),
      output(20) => mem_array(20)(360),
      output(21) => mem_array(21)(360),
      output(22) => mem_array(22)(360),
      output(23) => mem_array(23)(360),
      output(24) => mem_array(24)(360),
      output(25) => mem_array(25)(360),
      output(26) => mem_array(26)(360),
      output(27) => mem_array(27)(360),
      output(28) => mem_array(28)(360),
      output(29) => mem_array(29)(360),
      output(30) => mem_array(30)(360),
      output(31) => mem_array(31)(360),
      output(32) => mem_array(32)(360),
      output(33) => mem_array(33)(360),
      output(34) => mem_array(34)(360),
      output(35) => mem_array(35)(360)
      );
  rom361 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(361),
      output(0)  => mem_array(0)(361),
      output(1)  => mem_array(1)(361),
      output(2)  => mem_array(2)(361),
      output(3)  => mem_array(3)(361),
      output(4)  => mem_array(4)(361),
      output(5)  => mem_array(5)(361),
      output(6)  => mem_array(6)(361),
      output(7)  => mem_array(7)(361),
      output(8)  => mem_array(8)(361),
      output(9)  => mem_array(9)(361),
      output(10) => mem_array(10)(361),
      output(11) => mem_array(11)(361),
      output(12) => mem_array(12)(361),
      output(13) => mem_array(13)(361),
      output(14) => mem_array(14)(361),
      output(15) => mem_array(15)(361),
      output(16) => mem_array(16)(361),
      output(17) => mem_array(17)(361),
      output(18) => mem_array(18)(361),
      output(19) => mem_array(19)(361),
      output(20) => mem_array(20)(361),
      output(21) => mem_array(21)(361),
      output(22) => mem_array(22)(361),
      output(23) => mem_array(23)(361),
      output(24) => mem_array(24)(361),
      output(25) => mem_array(25)(361),
      output(26) => mem_array(26)(361),
      output(27) => mem_array(27)(361),
      output(28) => mem_array(28)(361),
      output(29) => mem_array(29)(361),
      output(30) => mem_array(30)(361),
      output(31) => mem_array(31)(361),
      output(32) => mem_array(32)(361),
      output(33) => mem_array(33)(361),
      output(34) => mem_array(34)(361),
      output(35) => mem_array(35)(361)
      );
  rom362 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(362),
      output(0)  => mem_array(0)(362),
      output(1)  => mem_array(1)(362),
      output(2)  => mem_array(2)(362),
      output(3)  => mem_array(3)(362),
      output(4)  => mem_array(4)(362),
      output(5)  => mem_array(5)(362),
      output(6)  => mem_array(6)(362),
      output(7)  => mem_array(7)(362),
      output(8)  => mem_array(8)(362),
      output(9)  => mem_array(9)(362),
      output(10) => mem_array(10)(362),
      output(11) => mem_array(11)(362),
      output(12) => mem_array(12)(362),
      output(13) => mem_array(13)(362),
      output(14) => mem_array(14)(362),
      output(15) => mem_array(15)(362),
      output(16) => mem_array(16)(362),
      output(17) => mem_array(17)(362),
      output(18) => mem_array(18)(362),
      output(19) => mem_array(19)(362),
      output(20) => mem_array(20)(362),
      output(21) => mem_array(21)(362),
      output(22) => mem_array(22)(362),
      output(23) => mem_array(23)(362),
      output(24) => mem_array(24)(362),
      output(25) => mem_array(25)(362),
      output(26) => mem_array(26)(362),
      output(27) => mem_array(27)(362),
      output(28) => mem_array(28)(362),
      output(29) => mem_array(29)(362),
      output(30) => mem_array(30)(362),
      output(31) => mem_array(31)(362),
      output(32) => mem_array(32)(362),
      output(33) => mem_array(33)(362),
      output(34) => mem_array(34)(362),
      output(35) => mem_array(35)(362)
      );
  rom363 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(363),
      output(0)  => mem_array(0)(363),
      output(1)  => mem_array(1)(363),
      output(2)  => mem_array(2)(363),
      output(3)  => mem_array(3)(363),
      output(4)  => mem_array(4)(363),
      output(5)  => mem_array(5)(363),
      output(6)  => mem_array(6)(363),
      output(7)  => mem_array(7)(363),
      output(8)  => mem_array(8)(363),
      output(9)  => mem_array(9)(363),
      output(10) => mem_array(10)(363),
      output(11) => mem_array(11)(363),
      output(12) => mem_array(12)(363),
      output(13) => mem_array(13)(363),
      output(14) => mem_array(14)(363),
      output(15) => mem_array(15)(363),
      output(16) => mem_array(16)(363),
      output(17) => mem_array(17)(363),
      output(18) => mem_array(18)(363),
      output(19) => mem_array(19)(363),
      output(20) => mem_array(20)(363),
      output(21) => mem_array(21)(363),
      output(22) => mem_array(22)(363),
      output(23) => mem_array(23)(363),
      output(24) => mem_array(24)(363),
      output(25) => mem_array(25)(363),
      output(26) => mem_array(26)(363),
      output(27) => mem_array(27)(363),
      output(28) => mem_array(28)(363),
      output(29) => mem_array(29)(363),
      output(30) => mem_array(30)(363),
      output(31) => mem_array(31)(363),
      output(32) => mem_array(32)(363),
      output(33) => mem_array(33)(363),
      output(34) => mem_array(34)(363),
      output(35) => mem_array(35)(363)
      );
  rom364 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(364),
      output(0)  => mem_array(0)(364),
      output(1)  => mem_array(1)(364),
      output(2)  => mem_array(2)(364),
      output(3)  => mem_array(3)(364),
      output(4)  => mem_array(4)(364),
      output(5)  => mem_array(5)(364),
      output(6)  => mem_array(6)(364),
      output(7)  => mem_array(7)(364),
      output(8)  => mem_array(8)(364),
      output(9)  => mem_array(9)(364),
      output(10) => mem_array(10)(364),
      output(11) => mem_array(11)(364),
      output(12) => mem_array(12)(364),
      output(13) => mem_array(13)(364),
      output(14) => mem_array(14)(364),
      output(15) => mem_array(15)(364),
      output(16) => mem_array(16)(364),
      output(17) => mem_array(17)(364),
      output(18) => mem_array(18)(364),
      output(19) => mem_array(19)(364),
      output(20) => mem_array(20)(364),
      output(21) => mem_array(21)(364),
      output(22) => mem_array(22)(364),
      output(23) => mem_array(23)(364),
      output(24) => mem_array(24)(364),
      output(25) => mem_array(25)(364),
      output(26) => mem_array(26)(364),
      output(27) => mem_array(27)(364),
      output(28) => mem_array(28)(364),
      output(29) => mem_array(29)(364),
      output(30) => mem_array(30)(364),
      output(31) => mem_array(31)(364),
      output(32) => mem_array(32)(364),
      output(33) => mem_array(33)(364),
      output(34) => mem_array(34)(364),
      output(35) => mem_array(35)(364)
      );
  rom365 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(365),
      output(0)  => mem_array(0)(365),
      output(1)  => mem_array(1)(365),
      output(2)  => mem_array(2)(365),
      output(3)  => mem_array(3)(365),
      output(4)  => mem_array(4)(365),
      output(5)  => mem_array(5)(365),
      output(6)  => mem_array(6)(365),
      output(7)  => mem_array(7)(365),
      output(8)  => mem_array(8)(365),
      output(9)  => mem_array(9)(365),
      output(10) => mem_array(10)(365),
      output(11) => mem_array(11)(365),
      output(12) => mem_array(12)(365),
      output(13) => mem_array(13)(365),
      output(14) => mem_array(14)(365),
      output(15) => mem_array(15)(365),
      output(16) => mem_array(16)(365),
      output(17) => mem_array(17)(365),
      output(18) => mem_array(18)(365),
      output(19) => mem_array(19)(365),
      output(20) => mem_array(20)(365),
      output(21) => mem_array(21)(365),
      output(22) => mem_array(22)(365),
      output(23) => mem_array(23)(365),
      output(24) => mem_array(24)(365),
      output(25) => mem_array(25)(365),
      output(26) => mem_array(26)(365),
      output(27) => mem_array(27)(365),
      output(28) => mem_array(28)(365),
      output(29) => mem_array(29)(365),
      output(30) => mem_array(30)(365),
      output(31) => mem_array(31)(365),
      output(32) => mem_array(32)(365),
      output(33) => mem_array(33)(365),
      output(34) => mem_array(34)(365),
      output(35) => mem_array(35)(365)
      );
  rom366 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(366),
      output(0)  => mem_array(0)(366),
      output(1)  => mem_array(1)(366),
      output(2)  => mem_array(2)(366),
      output(3)  => mem_array(3)(366),
      output(4)  => mem_array(4)(366),
      output(5)  => mem_array(5)(366),
      output(6)  => mem_array(6)(366),
      output(7)  => mem_array(7)(366),
      output(8)  => mem_array(8)(366),
      output(9)  => mem_array(9)(366),
      output(10) => mem_array(10)(366),
      output(11) => mem_array(11)(366),
      output(12) => mem_array(12)(366),
      output(13) => mem_array(13)(366),
      output(14) => mem_array(14)(366),
      output(15) => mem_array(15)(366),
      output(16) => mem_array(16)(366),
      output(17) => mem_array(17)(366),
      output(18) => mem_array(18)(366),
      output(19) => mem_array(19)(366),
      output(20) => mem_array(20)(366),
      output(21) => mem_array(21)(366),
      output(22) => mem_array(22)(366),
      output(23) => mem_array(23)(366),
      output(24) => mem_array(24)(366),
      output(25) => mem_array(25)(366),
      output(26) => mem_array(26)(366),
      output(27) => mem_array(27)(366),
      output(28) => mem_array(28)(366),
      output(29) => mem_array(29)(366),
      output(30) => mem_array(30)(366),
      output(31) => mem_array(31)(366),
      output(32) => mem_array(32)(366),
      output(33) => mem_array(33)(366),
      output(34) => mem_array(34)(366),
      output(35) => mem_array(35)(366)
      );
  rom367 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(367),
      output(0)  => mem_array(0)(367),
      output(1)  => mem_array(1)(367),
      output(2)  => mem_array(2)(367),
      output(3)  => mem_array(3)(367),
      output(4)  => mem_array(4)(367),
      output(5)  => mem_array(5)(367),
      output(6)  => mem_array(6)(367),
      output(7)  => mem_array(7)(367),
      output(8)  => mem_array(8)(367),
      output(9)  => mem_array(9)(367),
      output(10) => mem_array(10)(367),
      output(11) => mem_array(11)(367),
      output(12) => mem_array(12)(367),
      output(13) => mem_array(13)(367),
      output(14) => mem_array(14)(367),
      output(15) => mem_array(15)(367),
      output(16) => mem_array(16)(367),
      output(17) => mem_array(17)(367),
      output(18) => mem_array(18)(367),
      output(19) => mem_array(19)(367),
      output(20) => mem_array(20)(367),
      output(21) => mem_array(21)(367),
      output(22) => mem_array(22)(367),
      output(23) => mem_array(23)(367),
      output(24) => mem_array(24)(367),
      output(25) => mem_array(25)(367),
      output(26) => mem_array(26)(367),
      output(27) => mem_array(27)(367),
      output(28) => mem_array(28)(367),
      output(29) => mem_array(29)(367),
      output(30) => mem_array(30)(367),
      output(31) => mem_array(31)(367),
      output(32) => mem_array(32)(367),
      output(33) => mem_array(33)(367),
      output(34) => mem_array(34)(367),
      output(35) => mem_array(35)(367)
      );
  rom368 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(368),
      output(0)  => mem_array(0)(368),
      output(1)  => mem_array(1)(368),
      output(2)  => mem_array(2)(368),
      output(3)  => mem_array(3)(368),
      output(4)  => mem_array(4)(368),
      output(5)  => mem_array(5)(368),
      output(6)  => mem_array(6)(368),
      output(7)  => mem_array(7)(368),
      output(8)  => mem_array(8)(368),
      output(9)  => mem_array(9)(368),
      output(10) => mem_array(10)(368),
      output(11) => mem_array(11)(368),
      output(12) => mem_array(12)(368),
      output(13) => mem_array(13)(368),
      output(14) => mem_array(14)(368),
      output(15) => mem_array(15)(368),
      output(16) => mem_array(16)(368),
      output(17) => mem_array(17)(368),
      output(18) => mem_array(18)(368),
      output(19) => mem_array(19)(368),
      output(20) => mem_array(20)(368),
      output(21) => mem_array(21)(368),
      output(22) => mem_array(22)(368),
      output(23) => mem_array(23)(368),
      output(24) => mem_array(24)(368),
      output(25) => mem_array(25)(368),
      output(26) => mem_array(26)(368),
      output(27) => mem_array(27)(368),
      output(28) => mem_array(28)(368),
      output(29) => mem_array(29)(368),
      output(30) => mem_array(30)(368),
      output(31) => mem_array(31)(368),
      output(32) => mem_array(32)(368),
      output(33) => mem_array(33)(368),
      output(34) => mem_array(34)(368),
      output(35) => mem_array(35)(368)
      );
  rom369 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(369),
      output(0)  => mem_array(0)(369),
      output(1)  => mem_array(1)(369),
      output(2)  => mem_array(2)(369),
      output(3)  => mem_array(3)(369),
      output(4)  => mem_array(4)(369),
      output(5)  => mem_array(5)(369),
      output(6)  => mem_array(6)(369),
      output(7)  => mem_array(7)(369),
      output(8)  => mem_array(8)(369),
      output(9)  => mem_array(9)(369),
      output(10) => mem_array(10)(369),
      output(11) => mem_array(11)(369),
      output(12) => mem_array(12)(369),
      output(13) => mem_array(13)(369),
      output(14) => mem_array(14)(369),
      output(15) => mem_array(15)(369),
      output(16) => mem_array(16)(369),
      output(17) => mem_array(17)(369),
      output(18) => mem_array(18)(369),
      output(19) => mem_array(19)(369),
      output(20) => mem_array(20)(369),
      output(21) => mem_array(21)(369),
      output(22) => mem_array(22)(369),
      output(23) => mem_array(23)(369),
      output(24) => mem_array(24)(369),
      output(25) => mem_array(25)(369),
      output(26) => mem_array(26)(369),
      output(27) => mem_array(27)(369),
      output(28) => mem_array(28)(369),
      output(29) => mem_array(29)(369),
      output(30) => mem_array(30)(369),
      output(31) => mem_array(31)(369),
      output(32) => mem_array(32)(369),
      output(33) => mem_array(33)(369),
      output(34) => mem_array(34)(369),
      output(35) => mem_array(35)(369)
      );
  rom370 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(370),
      output(0)  => mem_array(0)(370),
      output(1)  => mem_array(1)(370),
      output(2)  => mem_array(2)(370),
      output(3)  => mem_array(3)(370),
      output(4)  => mem_array(4)(370),
      output(5)  => mem_array(5)(370),
      output(6)  => mem_array(6)(370),
      output(7)  => mem_array(7)(370),
      output(8)  => mem_array(8)(370),
      output(9)  => mem_array(9)(370),
      output(10) => mem_array(10)(370),
      output(11) => mem_array(11)(370),
      output(12) => mem_array(12)(370),
      output(13) => mem_array(13)(370),
      output(14) => mem_array(14)(370),
      output(15) => mem_array(15)(370),
      output(16) => mem_array(16)(370),
      output(17) => mem_array(17)(370),
      output(18) => mem_array(18)(370),
      output(19) => mem_array(19)(370),
      output(20) => mem_array(20)(370),
      output(21) => mem_array(21)(370),
      output(22) => mem_array(22)(370),
      output(23) => mem_array(23)(370),
      output(24) => mem_array(24)(370),
      output(25) => mem_array(25)(370),
      output(26) => mem_array(26)(370),
      output(27) => mem_array(27)(370),
      output(28) => mem_array(28)(370),
      output(29) => mem_array(29)(370),
      output(30) => mem_array(30)(370),
      output(31) => mem_array(31)(370),
      output(32) => mem_array(32)(370),
      output(33) => mem_array(33)(370),
      output(34) => mem_array(34)(370),
      output(35) => mem_array(35)(370)
      );
  rom371 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(371),
      output(0)  => mem_array(0)(371),
      output(1)  => mem_array(1)(371),
      output(2)  => mem_array(2)(371),
      output(3)  => mem_array(3)(371),
      output(4)  => mem_array(4)(371),
      output(5)  => mem_array(5)(371),
      output(6)  => mem_array(6)(371),
      output(7)  => mem_array(7)(371),
      output(8)  => mem_array(8)(371),
      output(9)  => mem_array(9)(371),
      output(10) => mem_array(10)(371),
      output(11) => mem_array(11)(371),
      output(12) => mem_array(12)(371),
      output(13) => mem_array(13)(371),
      output(14) => mem_array(14)(371),
      output(15) => mem_array(15)(371),
      output(16) => mem_array(16)(371),
      output(17) => mem_array(17)(371),
      output(18) => mem_array(18)(371),
      output(19) => mem_array(19)(371),
      output(20) => mem_array(20)(371),
      output(21) => mem_array(21)(371),
      output(22) => mem_array(22)(371),
      output(23) => mem_array(23)(371),
      output(24) => mem_array(24)(371),
      output(25) => mem_array(25)(371),
      output(26) => mem_array(26)(371),
      output(27) => mem_array(27)(371),
      output(28) => mem_array(28)(371),
      output(29) => mem_array(29)(371),
      output(30) => mem_array(30)(371),
      output(31) => mem_array(31)(371),
      output(32) => mem_array(32)(371),
      output(33) => mem_array(33)(371),
      output(34) => mem_array(34)(371),
      output(35) => mem_array(35)(371)
      );
  rom372 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(372),
      output(0)  => mem_array(0)(372),
      output(1)  => mem_array(1)(372),
      output(2)  => mem_array(2)(372),
      output(3)  => mem_array(3)(372),
      output(4)  => mem_array(4)(372),
      output(5)  => mem_array(5)(372),
      output(6)  => mem_array(6)(372),
      output(7)  => mem_array(7)(372),
      output(8)  => mem_array(8)(372),
      output(9)  => mem_array(9)(372),
      output(10) => mem_array(10)(372),
      output(11) => mem_array(11)(372),
      output(12) => mem_array(12)(372),
      output(13) => mem_array(13)(372),
      output(14) => mem_array(14)(372),
      output(15) => mem_array(15)(372),
      output(16) => mem_array(16)(372),
      output(17) => mem_array(17)(372),
      output(18) => mem_array(18)(372),
      output(19) => mem_array(19)(372),
      output(20) => mem_array(20)(372),
      output(21) => mem_array(21)(372),
      output(22) => mem_array(22)(372),
      output(23) => mem_array(23)(372),
      output(24) => mem_array(24)(372),
      output(25) => mem_array(25)(372),
      output(26) => mem_array(26)(372),
      output(27) => mem_array(27)(372),
      output(28) => mem_array(28)(372),
      output(29) => mem_array(29)(372),
      output(30) => mem_array(30)(372),
      output(31) => mem_array(31)(372),
      output(32) => mem_array(32)(372),
      output(33) => mem_array(33)(372),
      output(34) => mem_array(34)(372),
      output(35) => mem_array(35)(372)
      );
  rom373 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(373),
      output(0)  => mem_array(0)(373),
      output(1)  => mem_array(1)(373),
      output(2)  => mem_array(2)(373),
      output(3)  => mem_array(3)(373),
      output(4)  => mem_array(4)(373),
      output(5)  => mem_array(5)(373),
      output(6)  => mem_array(6)(373),
      output(7)  => mem_array(7)(373),
      output(8)  => mem_array(8)(373),
      output(9)  => mem_array(9)(373),
      output(10) => mem_array(10)(373),
      output(11) => mem_array(11)(373),
      output(12) => mem_array(12)(373),
      output(13) => mem_array(13)(373),
      output(14) => mem_array(14)(373),
      output(15) => mem_array(15)(373),
      output(16) => mem_array(16)(373),
      output(17) => mem_array(17)(373),
      output(18) => mem_array(18)(373),
      output(19) => mem_array(19)(373),
      output(20) => mem_array(20)(373),
      output(21) => mem_array(21)(373),
      output(22) => mem_array(22)(373),
      output(23) => mem_array(23)(373),
      output(24) => mem_array(24)(373),
      output(25) => mem_array(25)(373),
      output(26) => mem_array(26)(373),
      output(27) => mem_array(27)(373),
      output(28) => mem_array(28)(373),
      output(29) => mem_array(29)(373),
      output(30) => mem_array(30)(373),
      output(31) => mem_array(31)(373),
      output(32) => mem_array(32)(373),
      output(33) => mem_array(33)(373),
      output(34) => mem_array(34)(373),
      output(35) => mem_array(35)(373)
      );
  rom374 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(374),
      output(0)  => mem_array(0)(374),
      output(1)  => mem_array(1)(374),
      output(2)  => mem_array(2)(374),
      output(3)  => mem_array(3)(374),
      output(4)  => mem_array(4)(374),
      output(5)  => mem_array(5)(374),
      output(6)  => mem_array(6)(374),
      output(7)  => mem_array(7)(374),
      output(8)  => mem_array(8)(374),
      output(9)  => mem_array(9)(374),
      output(10) => mem_array(10)(374),
      output(11) => mem_array(11)(374),
      output(12) => mem_array(12)(374),
      output(13) => mem_array(13)(374),
      output(14) => mem_array(14)(374),
      output(15) => mem_array(15)(374),
      output(16) => mem_array(16)(374),
      output(17) => mem_array(17)(374),
      output(18) => mem_array(18)(374),
      output(19) => mem_array(19)(374),
      output(20) => mem_array(20)(374),
      output(21) => mem_array(21)(374),
      output(22) => mem_array(22)(374),
      output(23) => mem_array(23)(374),
      output(24) => mem_array(24)(374),
      output(25) => mem_array(25)(374),
      output(26) => mem_array(26)(374),
      output(27) => mem_array(27)(374),
      output(28) => mem_array(28)(374),
      output(29) => mem_array(29)(374),
      output(30) => mem_array(30)(374),
      output(31) => mem_array(31)(374),
      output(32) => mem_array(32)(374),
      output(33) => mem_array(33)(374),
      output(34) => mem_array(34)(374),
      output(35) => mem_array(35)(374)
      );
  rom375 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(375),
      output(0)  => mem_array(0)(375),
      output(1)  => mem_array(1)(375),
      output(2)  => mem_array(2)(375),
      output(3)  => mem_array(3)(375),
      output(4)  => mem_array(4)(375),
      output(5)  => mem_array(5)(375),
      output(6)  => mem_array(6)(375),
      output(7)  => mem_array(7)(375),
      output(8)  => mem_array(8)(375),
      output(9)  => mem_array(9)(375),
      output(10) => mem_array(10)(375),
      output(11) => mem_array(11)(375),
      output(12) => mem_array(12)(375),
      output(13) => mem_array(13)(375),
      output(14) => mem_array(14)(375),
      output(15) => mem_array(15)(375),
      output(16) => mem_array(16)(375),
      output(17) => mem_array(17)(375),
      output(18) => mem_array(18)(375),
      output(19) => mem_array(19)(375),
      output(20) => mem_array(20)(375),
      output(21) => mem_array(21)(375),
      output(22) => mem_array(22)(375),
      output(23) => mem_array(23)(375),
      output(24) => mem_array(24)(375),
      output(25) => mem_array(25)(375),
      output(26) => mem_array(26)(375),
      output(27) => mem_array(27)(375),
      output(28) => mem_array(28)(375),
      output(29) => mem_array(29)(375),
      output(30) => mem_array(30)(375),
      output(31) => mem_array(31)(375),
      output(32) => mem_array(32)(375),
      output(33) => mem_array(33)(375),
      output(34) => mem_array(34)(375),
      output(35) => mem_array(35)(375)
      );
  rom376 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(376),
      output(0)  => mem_array(0)(376),
      output(1)  => mem_array(1)(376),
      output(2)  => mem_array(2)(376),
      output(3)  => mem_array(3)(376),
      output(4)  => mem_array(4)(376),
      output(5)  => mem_array(5)(376),
      output(6)  => mem_array(6)(376),
      output(7)  => mem_array(7)(376),
      output(8)  => mem_array(8)(376),
      output(9)  => mem_array(9)(376),
      output(10) => mem_array(10)(376),
      output(11) => mem_array(11)(376),
      output(12) => mem_array(12)(376),
      output(13) => mem_array(13)(376),
      output(14) => mem_array(14)(376),
      output(15) => mem_array(15)(376),
      output(16) => mem_array(16)(376),
      output(17) => mem_array(17)(376),
      output(18) => mem_array(18)(376),
      output(19) => mem_array(19)(376),
      output(20) => mem_array(20)(376),
      output(21) => mem_array(21)(376),
      output(22) => mem_array(22)(376),
      output(23) => mem_array(23)(376),
      output(24) => mem_array(24)(376),
      output(25) => mem_array(25)(376),
      output(26) => mem_array(26)(376),
      output(27) => mem_array(27)(376),
      output(28) => mem_array(28)(376),
      output(29) => mem_array(29)(376),
      output(30) => mem_array(30)(376),
      output(31) => mem_array(31)(376),
      output(32) => mem_array(32)(376),
      output(33) => mem_array(33)(376),
      output(34) => mem_array(34)(376),
      output(35) => mem_array(35)(376)
      );
  rom377 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(377),
      output(0)  => mem_array(0)(377),
      output(1)  => mem_array(1)(377),
      output(2)  => mem_array(2)(377),
      output(3)  => mem_array(3)(377),
      output(4)  => mem_array(4)(377),
      output(5)  => mem_array(5)(377),
      output(6)  => mem_array(6)(377),
      output(7)  => mem_array(7)(377),
      output(8)  => mem_array(8)(377),
      output(9)  => mem_array(9)(377),
      output(10) => mem_array(10)(377),
      output(11) => mem_array(11)(377),
      output(12) => mem_array(12)(377),
      output(13) => mem_array(13)(377),
      output(14) => mem_array(14)(377),
      output(15) => mem_array(15)(377),
      output(16) => mem_array(16)(377),
      output(17) => mem_array(17)(377),
      output(18) => mem_array(18)(377),
      output(19) => mem_array(19)(377),
      output(20) => mem_array(20)(377),
      output(21) => mem_array(21)(377),
      output(22) => mem_array(22)(377),
      output(23) => mem_array(23)(377),
      output(24) => mem_array(24)(377),
      output(25) => mem_array(25)(377),
      output(26) => mem_array(26)(377),
      output(27) => mem_array(27)(377),
      output(28) => mem_array(28)(377),
      output(29) => mem_array(29)(377),
      output(30) => mem_array(30)(377),
      output(31) => mem_array(31)(377),
      output(32) => mem_array(32)(377),
      output(33) => mem_array(33)(377),
      output(34) => mem_array(34)(377),
      output(35) => mem_array(35)(377)
      );
  rom378 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(378),
      output(0)  => mem_array(0)(378),
      output(1)  => mem_array(1)(378),
      output(2)  => mem_array(2)(378),
      output(3)  => mem_array(3)(378),
      output(4)  => mem_array(4)(378),
      output(5)  => mem_array(5)(378),
      output(6)  => mem_array(6)(378),
      output(7)  => mem_array(7)(378),
      output(8)  => mem_array(8)(378),
      output(9)  => mem_array(9)(378),
      output(10) => mem_array(10)(378),
      output(11) => mem_array(11)(378),
      output(12) => mem_array(12)(378),
      output(13) => mem_array(13)(378),
      output(14) => mem_array(14)(378),
      output(15) => mem_array(15)(378),
      output(16) => mem_array(16)(378),
      output(17) => mem_array(17)(378),
      output(18) => mem_array(18)(378),
      output(19) => mem_array(19)(378),
      output(20) => mem_array(20)(378),
      output(21) => mem_array(21)(378),
      output(22) => mem_array(22)(378),
      output(23) => mem_array(23)(378),
      output(24) => mem_array(24)(378),
      output(25) => mem_array(25)(378),
      output(26) => mem_array(26)(378),
      output(27) => mem_array(27)(378),
      output(28) => mem_array(28)(378),
      output(29) => mem_array(29)(378),
      output(30) => mem_array(30)(378),
      output(31) => mem_array(31)(378),
      output(32) => mem_array(32)(378),
      output(33) => mem_array(33)(378),
      output(34) => mem_array(34)(378),
      output(35) => mem_array(35)(378)
      );
  rom379 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(379),
      output(0)  => mem_array(0)(379),
      output(1)  => mem_array(1)(379),
      output(2)  => mem_array(2)(379),
      output(3)  => mem_array(3)(379),
      output(4)  => mem_array(4)(379),
      output(5)  => mem_array(5)(379),
      output(6)  => mem_array(6)(379),
      output(7)  => mem_array(7)(379),
      output(8)  => mem_array(8)(379),
      output(9)  => mem_array(9)(379),
      output(10) => mem_array(10)(379),
      output(11) => mem_array(11)(379),
      output(12) => mem_array(12)(379),
      output(13) => mem_array(13)(379),
      output(14) => mem_array(14)(379),
      output(15) => mem_array(15)(379),
      output(16) => mem_array(16)(379),
      output(17) => mem_array(17)(379),
      output(18) => mem_array(18)(379),
      output(19) => mem_array(19)(379),
      output(20) => mem_array(20)(379),
      output(21) => mem_array(21)(379),
      output(22) => mem_array(22)(379),
      output(23) => mem_array(23)(379),
      output(24) => mem_array(24)(379),
      output(25) => mem_array(25)(379),
      output(26) => mem_array(26)(379),
      output(27) => mem_array(27)(379),
      output(28) => mem_array(28)(379),
      output(29) => mem_array(29)(379),
      output(30) => mem_array(30)(379),
      output(31) => mem_array(31)(379),
      output(32) => mem_array(32)(379),
      output(33) => mem_array(33)(379),
      output(34) => mem_array(34)(379),
      output(35) => mem_array(35)(379)
      );
  rom380 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(380),
      output(0)  => mem_array(0)(380),
      output(1)  => mem_array(1)(380),
      output(2)  => mem_array(2)(380),
      output(3)  => mem_array(3)(380),
      output(4)  => mem_array(4)(380),
      output(5)  => mem_array(5)(380),
      output(6)  => mem_array(6)(380),
      output(7)  => mem_array(7)(380),
      output(8)  => mem_array(8)(380),
      output(9)  => mem_array(9)(380),
      output(10) => mem_array(10)(380),
      output(11) => mem_array(11)(380),
      output(12) => mem_array(12)(380),
      output(13) => mem_array(13)(380),
      output(14) => mem_array(14)(380),
      output(15) => mem_array(15)(380),
      output(16) => mem_array(16)(380),
      output(17) => mem_array(17)(380),
      output(18) => mem_array(18)(380),
      output(19) => mem_array(19)(380),
      output(20) => mem_array(20)(380),
      output(21) => mem_array(21)(380),
      output(22) => mem_array(22)(380),
      output(23) => mem_array(23)(380),
      output(24) => mem_array(24)(380),
      output(25) => mem_array(25)(380),
      output(26) => mem_array(26)(380),
      output(27) => mem_array(27)(380),
      output(28) => mem_array(28)(380),
      output(29) => mem_array(29)(380),
      output(30) => mem_array(30)(380),
      output(31) => mem_array(31)(380),
      output(32) => mem_array(32)(380),
      output(33) => mem_array(33)(380),
      output(34) => mem_array(34)(380),
      output(35) => mem_array(35)(380)
      );
  rom381 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(381),
      output(0)  => mem_array(0)(381),
      output(1)  => mem_array(1)(381),
      output(2)  => mem_array(2)(381),
      output(3)  => mem_array(3)(381),
      output(4)  => mem_array(4)(381),
      output(5)  => mem_array(5)(381),
      output(6)  => mem_array(6)(381),
      output(7)  => mem_array(7)(381),
      output(8)  => mem_array(8)(381),
      output(9)  => mem_array(9)(381),
      output(10) => mem_array(10)(381),
      output(11) => mem_array(11)(381),
      output(12) => mem_array(12)(381),
      output(13) => mem_array(13)(381),
      output(14) => mem_array(14)(381),
      output(15) => mem_array(15)(381),
      output(16) => mem_array(16)(381),
      output(17) => mem_array(17)(381),
      output(18) => mem_array(18)(381),
      output(19) => mem_array(19)(381),
      output(20) => mem_array(20)(381),
      output(21) => mem_array(21)(381),
      output(22) => mem_array(22)(381),
      output(23) => mem_array(23)(381),
      output(24) => mem_array(24)(381),
      output(25) => mem_array(25)(381),
      output(26) => mem_array(26)(381),
      output(27) => mem_array(27)(381),
      output(28) => mem_array(28)(381),
      output(29) => mem_array(29)(381),
      output(30) => mem_array(30)(381),
      output(31) => mem_array(31)(381),
      output(32) => mem_array(32)(381),
      output(33) => mem_array(33)(381),
      output(34) => mem_array(34)(381),
      output(35) => mem_array(35)(381)
      );
  rom382 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(382),
      output(0)  => mem_array(0)(382),
      output(1)  => mem_array(1)(382),
      output(2)  => mem_array(2)(382),
      output(3)  => mem_array(3)(382),
      output(4)  => mem_array(4)(382),
      output(5)  => mem_array(5)(382),
      output(6)  => mem_array(6)(382),
      output(7)  => mem_array(7)(382),
      output(8)  => mem_array(8)(382),
      output(9)  => mem_array(9)(382),
      output(10) => mem_array(10)(382),
      output(11) => mem_array(11)(382),
      output(12) => mem_array(12)(382),
      output(13) => mem_array(13)(382),
      output(14) => mem_array(14)(382),
      output(15) => mem_array(15)(382),
      output(16) => mem_array(16)(382),
      output(17) => mem_array(17)(382),
      output(18) => mem_array(18)(382),
      output(19) => mem_array(19)(382),
      output(20) => mem_array(20)(382),
      output(21) => mem_array(21)(382),
      output(22) => mem_array(22)(382),
      output(23) => mem_array(23)(382),
      output(24) => mem_array(24)(382),
      output(25) => mem_array(25)(382),
      output(26) => mem_array(26)(382),
      output(27) => mem_array(27)(382),
      output(28) => mem_array(28)(382),
      output(29) => mem_array(29)(382),
      output(30) => mem_array(30)(382),
      output(31) => mem_array(31)(382),
      output(32) => mem_array(32)(382),
      output(33) => mem_array(33)(382),
      output(34) => mem_array(34)(382),
      output(35) => mem_array(35)(382)
      );
  rom383 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(383),
      output(0)  => mem_array(0)(383),
      output(1)  => mem_array(1)(383),
      output(2)  => mem_array(2)(383),
      output(3)  => mem_array(3)(383),
      output(4)  => mem_array(4)(383),
      output(5)  => mem_array(5)(383),
      output(6)  => mem_array(6)(383),
      output(7)  => mem_array(7)(383),
      output(8)  => mem_array(8)(383),
      output(9)  => mem_array(9)(383),
      output(10) => mem_array(10)(383),
      output(11) => mem_array(11)(383),
      output(12) => mem_array(12)(383),
      output(13) => mem_array(13)(383),
      output(14) => mem_array(14)(383),
      output(15) => mem_array(15)(383),
      output(16) => mem_array(16)(383),
      output(17) => mem_array(17)(383),
      output(18) => mem_array(18)(383),
      output(19) => mem_array(19)(383),
      output(20) => mem_array(20)(383),
      output(21) => mem_array(21)(383),
      output(22) => mem_array(22)(383),
      output(23) => mem_array(23)(383),
      output(24) => mem_array(24)(383),
      output(25) => mem_array(25)(383),
      output(26) => mem_array(26)(383),
      output(27) => mem_array(27)(383),
      output(28) => mem_array(28)(383),
      output(29) => mem_array(29)(383),
      output(30) => mem_array(30)(383),
      output(31) => mem_array(31)(383),
      output(32) => mem_array(32)(383),
      output(33) => mem_array(33)(383),
      output(34) => mem_array(34)(383),
      output(35) => mem_array(35)(383)
      );
  rom384 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(384),
      output(0)  => mem_array(0)(384),
      output(1)  => mem_array(1)(384),
      output(2)  => mem_array(2)(384),
      output(3)  => mem_array(3)(384),
      output(4)  => mem_array(4)(384),
      output(5)  => mem_array(5)(384),
      output(6)  => mem_array(6)(384),
      output(7)  => mem_array(7)(384),
      output(8)  => mem_array(8)(384),
      output(9)  => mem_array(9)(384),
      output(10) => mem_array(10)(384),
      output(11) => mem_array(11)(384),
      output(12) => mem_array(12)(384),
      output(13) => mem_array(13)(384),
      output(14) => mem_array(14)(384),
      output(15) => mem_array(15)(384),
      output(16) => mem_array(16)(384),
      output(17) => mem_array(17)(384),
      output(18) => mem_array(18)(384),
      output(19) => mem_array(19)(384),
      output(20) => mem_array(20)(384),
      output(21) => mem_array(21)(384),
      output(22) => mem_array(22)(384),
      output(23) => mem_array(23)(384),
      output(24) => mem_array(24)(384),
      output(25) => mem_array(25)(384),
      output(26) => mem_array(26)(384),
      output(27) => mem_array(27)(384),
      output(28) => mem_array(28)(384),
      output(29) => mem_array(29)(384),
      output(30) => mem_array(30)(384),
      output(31) => mem_array(31)(384),
      output(32) => mem_array(32)(384),
      output(33) => mem_array(33)(384),
      output(34) => mem_array(34)(384),
      output(35) => mem_array(35)(384)
      );
  rom385 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(385),
      output(0)  => mem_array(0)(385),
      output(1)  => mem_array(1)(385),
      output(2)  => mem_array(2)(385),
      output(3)  => mem_array(3)(385),
      output(4)  => mem_array(4)(385),
      output(5)  => mem_array(5)(385),
      output(6)  => mem_array(6)(385),
      output(7)  => mem_array(7)(385),
      output(8)  => mem_array(8)(385),
      output(9)  => mem_array(9)(385),
      output(10) => mem_array(10)(385),
      output(11) => mem_array(11)(385),
      output(12) => mem_array(12)(385),
      output(13) => mem_array(13)(385),
      output(14) => mem_array(14)(385),
      output(15) => mem_array(15)(385),
      output(16) => mem_array(16)(385),
      output(17) => mem_array(17)(385),
      output(18) => mem_array(18)(385),
      output(19) => mem_array(19)(385),
      output(20) => mem_array(20)(385),
      output(21) => mem_array(21)(385),
      output(22) => mem_array(22)(385),
      output(23) => mem_array(23)(385),
      output(24) => mem_array(24)(385),
      output(25) => mem_array(25)(385),
      output(26) => mem_array(26)(385),
      output(27) => mem_array(27)(385),
      output(28) => mem_array(28)(385),
      output(29) => mem_array(29)(385),
      output(30) => mem_array(30)(385),
      output(31) => mem_array(31)(385),
      output(32) => mem_array(32)(385),
      output(33) => mem_array(33)(385),
      output(34) => mem_array(34)(385),
      output(35) => mem_array(35)(385)
      );
  rom386 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(386),
      output(0)  => mem_array(0)(386),
      output(1)  => mem_array(1)(386),
      output(2)  => mem_array(2)(386),
      output(3)  => mem_array(3)(386),
      output(4)  => mem_array(4)(386),
      output(5)  => mem_array(5)(386),
      output(6)  => mem_array(6)(386),
      output(7)  => mem_array(7)(386),
      output(8)  => mem_array(8)(386),
      output(9)  => mem_array(9)(386),
      output(10) => mem_array(10)(386),
      output(11) => mem_array(11)(386),
      output(12) => mem_array(12)(386),
      output(13) => mem_array(13)(386),
      output(14) => mem_array(14)(386),
      output(15) => mem_array(15)(386),
      output(16) => mem_array(16)(386),
      output(17) => mem_array(17)(386),
      output(18) => mem_array(18)(386),
      output(19) => mem_array(19)(386),
      output(20) => mem_array(20)(386),
      output(21) => mem_array(21)(386),
      output(22) => mem_array(22)(386),
      output(23) => mem_array(23)(386),
      output(24) => mem_array(24)(386),
      output(25) => mem_array(25)(386),
      output(26) => mem_array(26)(386),
      output(27) => mem_array(27)(386),
      output(28) => mem_array(28)(386),
      output(29) => mem_array(29)(386),
      output(30) => mem_array(30)(386),
      output(31) => mem_array(31)(386),
      output(32) => mem_array(32)(386),
      output(33) => mem_array(33)(386),
      output(34) => mem_array(34)(386),
      output(35) => mem_array(35)(386)
      );
  rom387 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(387),
      output(0)  => mem_array(0)(387),
      output(1)  => mem_array(1)(387),
      output(2)  => mem_array(2)(387),
      output(3)  => mem_array(3)(387),
      output(4)  => mem_array(4)(387),
      output(5)  => mem_array(5)(387),
      output(6)  => mem_array(6)(387),
      output(7)  => mem_array(7)(387),
      output(8)  => mem_array(8)(387),
      output(9)  => mem_array(9)(387),
      output(10) => mem_array(10)(387),
      output(11) => mem_array(11)(387),
      output(12) => mem_array(12)(387),
      output(13) => mem_array(13)(387),
      output(14) => mem_array(14)(387),
      output(15) => mem_array(15)(387),
      output(16) => mem_array(16)(387),
      output(17) => mem_array(17)(387),
      output(18) => mem_array(18)(387),
      output(19) => mem_array(19)(387),
      output(20) => mem_array(20)(387),
      output(21) => mem_array(21)(387),
      output(22) => mem_array(22)(387),
      output(23) => mem_array(23)(387),
      output(24) => mem_array(24)(387),
      output(25) => mem_array(25)(387),
      output(26) => mem_array(26)(387),
      output(27) => mem_array(27)(387),
      output(28) => mem_array(28)(387),
      output(29) => mem_array(29)(387),
      output(30) => mem_array(30)(387),
      output(31) => mem_array(31)(387),
      output(32) => mem_array(32)(387),
      output(33) => mem_array(33)(387),
      output(34) => mem_array(34)(387),
      output(35) => mem_array(35)(387)
      );
  rom388 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(388),
      output(0)  => mem_array(0)(388),
      output(1)  => mem_array(1)(388),
      output(2)  => mem_array(2)(388),
      output(3)  => mem_array(3)(388),
      output(4)  => mem_array(4)(388),
      output(5)  => mem_array(5)(388),
      output(6)  => mem_array(6)(388),
      output(7)  => mem_array(7)(388),
      output(8)  => mem_array(8)(388),
      output(9)  => mem_array(9)(388),
      output(10) => mem_array(10)(388),
      output(11) => mem_array(11)(388),
      output(12) => mem_array(12)(388),
      output(13) => mem_array(13)(388),
      output(14) => mem_array(14)(388),
      output(15) => mem_array(15)(388),
      output(16) => mem_array(16)(388),
      output(17) => mem_array(17)(388),
      output(18) => mem_array(18)(388),
      output(19) => mem_array(19)(388),
      output(20) => mem_array(20)(388),
      output(21) => mem_array(21)(388),
      output(22) => mem_array(22)(388),
      output(23) => mem_array(23)(388),
      output(24) => mem_array(24)(388),
      output(25) => mem_array(25)(388),
      output(26) => mem_array(26)(388),
      output(27) => mem_array(27)(388),
      output(28) => mem_array(28)(388),
      output(29) => mem_array(29)(388),
      output(30) => mem_array(30)(388),
      output(31) => mem_array(31)(388),
      output(32) => mem_array(32)(388),
      output(33) => mem_array(33)(388),
      output(34) => mem_array(34)(388),
      output(35) => mem_array(35)(388)
      );
  rom389 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(389),
      output(0)  => mem_array(0)(389),
      output(1)  => mem_array(1)(389),
      output(2)  => mem_array(2)(389),
      output(3)  => mem_array(3)(389),
      output(4)  => mem_array(4)(389),
      output(5)  => mem_array(5)(389),
      output(6)  => mem_array(6)(389),
      output(7)  => mem_array(7)(389),
      output(8)  => mem_array(8)(389),
      output(9)  => mem_array(9)(389),
      output(10) => mem_array(10)(389),
      output(11) => mem_array(11)(389),
      output(12) => mem_array(12)(389),
      output(13) => mem_array(13)(389),
      output(14) => mem_array(14)(389),
      output(15) => mem_array(15)(389),
      output(16) => mem_array(16)(389),
      output(17) => mem_array(17)(389),
      output(18) => mem_array(18)(389),
      output(19) => mem_array(19)(389),
      output(20) => mem_array(20)(389),
      output(21) => mem_array(21)(389),
      output(22) => mem_array(22)(389),
      output(23) => mem_array(23)(389),
      output(24) => mem_array(24)(389),
      output(25) => mem_array(25)(389),
      output(26) => mem_array(26)(389),
      output(27) => mem_array(27)(389),
      output(28) => mem_array(28)(389),
      output(29) => mem_array(29)(389),
      output(30) => mem_array(30)(389),
      output(31) => mem_array(31)(389),
      output(32) => mem_array(32)(389),
      output(33) => mem_array(33)(389),
      output(34) => mem_array(34)(389),
      output(35) => mem_array(35)(389)
      );
  rom390 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(390),
      output(0)  => mem_array(0)(390),
      output(1)  => mem_array(1)(390),
      output(2)  => mem_array(2)(390),
      output(3)  => mem_array(3)(390),
      output(4)  => mem_array(4)(390),
      output(5)  => mem_array(5)(390),
      output(6)  => mem_array(6)(390),
      output(7)  => mem_array(7)(390),
      output(8)  => mem_array(8)(390),
      output(9)  => mem_array(9)(390),
      output(10) => mem_array(10)(390),
      output(11) => mem_array(11)(390),
      output(12) => mem_array(12)(390),
      output(13) => mem_array(13)(390),
      output(14) => mem_array(14)(390),
      output(15) => mem_array(15)(390),
      output(16) => mem_array(16)(390),
      output(17) => mem_array(17)(390),
      output(18) => mem_array(18)(390),
      output(19) => mem_array(19)(390),
      output(20) => mem_array(20)(390),
      output(21) => mem_array(21)(390),
      output(22) => mem_array(22)(390),
      output(23) => mem_array(23)(390),
      output(24) => mem_array(24)(390),
      output(25) => mem_array(25)(390),
      output(26) => mem_array(26)(390),
      output(27) => mem_array(27)(390),
      output(28) => mem_array(28)(390),
      output(29) => mem_array(29)(390),
      output(30) => mem_array(30)(390),
      output(31) => mem_array(31)(390),
      output(32) => mem_array(32)(390),
      output(33) => mem_array(33)(390),
      output(34) => mem_array(34)(390),
      output(35) => mem_array(35)(390)
      );
  rom391 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(391),
      output(0)  => mem_array(0)(391),
      output(1)  => mem_array(1)(391),
      output(2)  => mem_array(2)(391),
      output(3)  => mem_array(3)(391),
      output(4)  => mem_array(4)(391),
      output(5)  => mem_array(5)(391),
      output(6)  => mem_array(6)(391),
      output(7)  => mem_array(7)(391),
      output(8)  => mem_array(8)(391),
      output(9)  => mem_array(9)(391),
      output(10) => mem_array(10)(391),
      output(11) => mem_array(11)(391),
      output(12) => mem_array(12)(391),
      output(13) => mem_array(13)(391),
      output(14) => mem_array(14)(391),
      output(15) => mem_array(15)(391),
      output(16) => mem_array(16)(391),
      output(17) => mem_array(17)(391),
      output(18) => mem_array(18)(391),
      output(19) => mem_array(19)(391),
      output(20) => mem_array(20)(391),
      output(21) => mem_array(21)(391),
      output(22) => mem_array(22)(391),
      output(23) => mem_array(23)(391),
      output(24) => mem_array(24)(391),
      output(25) => mem_array(25)(391),
      output(26) => mem_array(26)(391),
      output(27) => mem_array(27)(391),
      output(28) => mem_array(28)(391),
      output(29) => mem_array(29)(391),
      output(30) => mem_array(30)(391),
      output(31) => mem_array(31)(391),
      output(32) => mem_array(32)(391),
      output(33) => mem_array(33)(391),
      output(34) => mem_array(34)(391),
      output(35) => mem_array(35)(391)
      );
  rom392 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(392),
      output(0)  => mem_array(0)(392),
      output(1)  => mem_array(1)(392),
      output(2)  => mem_array(2)(392),
      output(3)  => mem_array(3)(392),
      output(4)  => mem_array(4)(392),
      output(5)  => mem_array(5)(392),
      output(6)  => mem_array(6)(392),
      output(7)  => mem_array(7)(392),
      output(8)  => mem_array(8)(392),
      output(9)  => mem_array(9)(392),
      output(10) => mem_array(10)(392),
      output(11) => mem_array(11)(392),
      output(12) => mem_array(12)(392),
      output(13) => mem_array(13)(392),
      output(14) => mem_array(14)(392),
      output(15) => mem_array(15)(392),
      output(16) => mem_array(16)(392),
      output(17) => mem_array(17)(392),
      output(18) => mem_array(18)(392),
      output(19) => mem_array(19)(392),
      output(20) => mem_array(20)(392),
      output(21) => mem_array(21)(392),
      output(22) => mem_array(22)(392),
      output(23) => mem_array(23)(392),
      output(24) => mem_array(24)(392),
      output(25) => mem_array(25)(392),
      output(26) => mem_array(26)(392),
      output(27) => mem_array(27)(392),
      output(28) => mem_array(28)(392),
      output(29) => mem_array(29)(392),
      output(30) => mem_array(30)(392),
      output(31) => mem_array(31)(392),
      output(32) => mem_array(32)(392),
      output(33) => mem_array(33)(392),
      output(34) => mem_array(34)(392),
      output(35) => mem_array(35)(392)
      );
  rom393 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(393),
      output(0)  => mem_array(0)(393),
      output(1)  => mem_array(1)(393),
      output(2)  => mem_array(2)(393),
      output(3)  => mem_array(3)(393),
      output(4)  => mem_array(4)(393),
      output(5)  => mem_array(5)(393),
      output(6)  => mem_array(6)(393),
      output(7)  => mem_array(7)(393),
      output(8)  => mem_array(8)(393),
      output(9)  => mem_array(9)(393),
      output(10) => mem_array(10)(393),
      output(11) => mem_array(11)(393),
      output(12) => mem_array(12)(393),
      output(13) => mem_array(13)(393),
      output(14) => mem_array(14)(393),
      output(15) => mem_array(15)(393),
      output(16) => mem_array(16)(393),
      output(17) => mem_array(17)(393),
      output(18) => mem_array(18)(393),
      output(19) => mem_array(19)(393),
      output(20) => mem_array(20)(393),
      output(21) => mem_array(21)(393),
      output(22) => mem_array(22)(393),
      output(23) => mem_array(23)(393),
      output(24) => mem_array(24)(393),
      output(25) => mem_array(25)(393),
      output(26) => mem_array(26)(393),
      output(27) => mem_array(27)(393),
      output(28) => mem_array(28)(393),
      output(29) => mem_array(29)(393),
      output(30) => mem_array(30)(393),
      output(31) => mem_array(31)(393),
      output(32) => mem_array(32)(393),
      output(33) => mem_array(33)(393),
      output(34) => mem_array(34)(393),
      output(35) => mem_array(35)(393)
      );
  rom394 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(394),
      output(0)  => mem_array(0)(394),
      output(1)  => mem_array(1)(394),
      output(2)  => mem_array(2)(394),
      output(3)  => mem_array(3)(394),
      output(4)  => mem_array(4)(394),
      output(5)  => mem_array(5)(394),
      output(6)  => mem_array(6)(394),
      output(7)  => mem_array(7)(394),
      output(8)  => mem_array(8)(394),
      output(9)  => mem_array(9)(394),
      output(10) => mem_array(10)(394),
      output(11) => mem_array(11)(394),
      output(12) => mem_array(12)(394),
      output(13) => mem_array(13)(394),
      output(14) => mem_array(14)(394),
      output(15) => mem_array(15)(394),
      output(16) => mem_array(16)(394),
      output(17) => mem_array(17)(394),
      output(18) => mem_array(18)(394),
      output(19) => mem_array(19)(394),
      output(20) => mem_array(20)(394),
      output(21) => mem_array(21)(394),
      output(22) => mem_array(22)(394),
      output(23) => mem_array(23)(394),
      output(24) => mem_array(24)(394),
      output(25) => mem_array(25)(394),
      output(26) => mem_array(26)(394),
      output(27) => mem_array(27)(394),
      output(28) => mem_array(28)(394),
      output(29) => mem_array(29)(394),
      output(30) => mem_array(30)(394),
      output(31) => mem_array(31)(394),
      output(32) => mem_array(32)(394),
      output(33) => mem_array(33)(394),
      output(34) => mem_array(34)(394),
      output(35) => mem_array(35)(394)
      );
  rom395 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(395),
      output(0)  => mem_array(0)(395),
      output(1)  => mem_array(1)(395),
      output(2)  => mem_array(2)(395),
      output(3)  => mem_array(3)(395),
      output(4)  => mem_array(4)(395),
      output(5)  => mem_array(5)(395),
      output(6)  => mem_array(6)(395),
      output(7)  => mem_array(7)(395),
      output(8)  => mem_array(8)(395),
      output(9)  => mem_array(9)(395),
      output(10) => mem_array(10)(395),
      output(11) => mem_array(11)(395),
      output(12) => mem_array(12)(395),
      output(13) => mem_array(13)(395),
      output(14) => mem_array(14)(395),
      output(15) => mem_array(15)(395),
      output(16) => mem_array(16)(395),
      output(17) => mem_array(17)(395),
      output(18) => mem_array(18)(395),
      output(19) => mem_array(19)(395),
      output(20) => mem_array(20)(395),
      output(21) => mem_array(21)(395),
      output(22) => mem_array(22)(395),
      output(23) => mem_array(23)(395),
      output(24) => mem_array(24)(395),
      output(25) => mem_array(25)(395),
      output(26) => mem_array(26)(395),
      output(27) => mem_array(27)(395),
      output(28) => mem_array(28)(395),
      output(29) => mem_array(29)(395),
      output(30) => mem_array(30)(395),
      output(31) => mem_array(31)(395),
      output(32) => mem_array(32)(395),
      output(33) => mem_array(33)(395),
      output(34) => mem_array(34)(395),
      output(35) => mem_array(35)(395)
      );
  rom396 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(396),
      output(0)  => mem_array(0)(396),
      output(1)  => mem_array(1)(396),
      output(2)  => mem_array(2)(396),
      output(3)  => mem_array(3)(396),
      output(4)  => mem_array(4)(396),
      output(5)  => mem_array(5)(396),
      output(6)  => mem_array(6)(396),
      output(7)  => mem_array(7)(396),
      output(8)  => mem_array(8)(396),
      output(9)  => mem_array(9)(396),
      output(10) => mem_array(10)(396),
      output(11) => mem_array(11)(396),
      output(12) => mem_array(12)(396),
      output(13) => mem_array(13)(396),
      output(14) => mem_array(14)(396),
      output(15) => mem_array(15)(396),
      output(16) => mem_array(16)(396),
      output(17) => mem_array(17)(396),
      output(18) => mem_array(18)(396),
      output(19) => mem_array(19)(396),
      output(20) => mem_array(20)(396),
      output(21) => mem_array(21)(396),
      output(22) => mem_array(22)(396),
      output(23) => mem_array(23)(396),
      output(24) => mem_array(24)(396),
      output(25) => mem_array(25)(396),
      output(26) => mem_array(26)(396),
      output(27) => mem_array(27)(396),
      output(28) => mem_array(28)(396),
      output(29) => mem_array(29)(396),
      output(30) => mem_array(30)(396),
      output(31) => mem_array(31)(396),
      output(32) => mem_array(32)(396),
      output(33) => mem_array(33)(396),
      output(34) => mem_array(34)(396),
      output(35) => mem_array(35)(396)
      );
  rom397 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(397),
      output(0)  => mem_array(0)(397),
      output(1)  => mem_array(1)(397),
      output(2)  => mem_array(2)(397),
      output(3)  => mem_array(3)(397),
      output(4)  => mem_array(4)(397),
      output(5)  => mem_array(5)(397),
      output(6)  => mem_array(6)(397),
      output(7)  => mem_array(7)(397),
      output(8)  => mem_array(8)(397),
      output(9)  => mem_array(9)(397),
      output(10) => mem_array(10)(397),
      output(11) => mem_array(11)(397),
      output(12) => mem_array(12)(397),
      output(13) => mem_array(13)(397),
      output(14) => mem_array(14)(397),
      output(15) => mem_array(15)(397),
      output(16) => mem_array(16)(397),
      output(17) => mem_array(17)(397),
      output(18) => mem_array(18)(397),
      output(19) => mem_array(19)(397),
      output(20) => mem_array(20)(397),
      output(21) => mem_array(21)(397),
      output(22) => mem_array(22)(397),
      output(23) => mem_array(23)(397),
      output(24) => mem_array(24)(397),
      output(25) => mem_array(25)(397),
      output(26) => mem_array(26)(397),
      output(27) => mem_array(27)(397),
      output(28) => mem_array(28)(397),
      output(29) => mem_array(29)(397),
      output(30) => mem_array(30)(397),
      output(31) => mem_array(31)(397),
      output(32) => mem_array(32)(397),
      output(33) => mem_array(33)(397),
      output(34) => mem_array(34)(397),
      output(35) => mem_array(35)(397)
      );
  rom398 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(398),
      output(0)  => mem_array(0)(398),
      output(1)  => mem_array(1)(398),
      output(2)  => mem_array(2)(398),
      output(3)  => mem_array(3)(398),
      output(4)  => mem_array(4)(398),
      output(5)  => mem_array(5)(398),
      output(6)  => mem_array(6)(398),
      output(7)  => mem_array(7)(398),
      output(8)  => mem_array(8)(398),
      output(9)  => mem_array(9)(398),
      output(10) => mem_array(10)(398),
      output(11) => mem_array(11)(398),
      output(12) => mem_array(12)(398),
      output(13) => mem_array(13)(398),
      output(14) => mem_array(14)(398),
      output(15) => mem_array(15)(398),
      output(16) => mem_array(16)(398),
      output(17) => mem_array(17)(398),
      output(18) => mem_array(18)(398),
      output(19) => mem_array(19)(398),
      output(20) => mem_array(20)(398),
      output(21) => mem_array(21)(398),
      output(22) => mem_array(22)(398),
      output(23) => mem_array(23)(398),
      output(24) => mem_array(24)(398),
      output(25) => mem_array(25)(398),
      output(26) => mem_array(26)(398),
      output(27) => mem_array(27)(398),
      output(28) => mem_array(28)(398),
      output(29) => mem_array(29)(398),
      output(30) => mem_array(30)(398),
      output(31) => mem_array(31)(398),
      output(32) => mem_array(32)(398),
      output(33) => mem_array(33)(398),
      output(34) => mem_array(34)(398),
      output(35) => mem_array(35)(398)
      );
  rom399 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(399),
      output(0)  => mem_array(0)(399),
      output(1)  => mem_array(1)(399),
      output(2)  => mem_array(2)(399),
      output(3)  => mem_array(3)(399),
      output(4)  => mem_array(4)(399),
      output(5)  => mem_array(5)(399),
      output(6)  => mem_array(6)(399),
      output(7)  => mem_array(7)(399),
      output(8)  => mem_array(8)(399),
      output(9)  => mem_array(9)(399),
      output(10) => mem_array(10)(399),
      output(11) => mem_array(11)(399),
      output(12) => mem_array(12)(399),
      output(13) => mem_array(13)(399),
      output(14) => mem_array(14)(399),
      output(15) => mem_array(15)(399),
      output(16) => mem_array(16)(399),
      output(17) => mem_array(17)(399),
      output(18) => mem_array(18)(399),
      output(19) => mem_array(19)(399),
      output(20) => mem_array(20)(399),
      output(21) => mem_array(21)(399),
      output(22) => mem_array(22)(399),
      output(23) => mem_array(23)(399),
      output(24) => mem_array(24)(399),
      output(25) => mem_array(25)(399),
      output(26) => mem_array(26)(399),
      output(27) => mem_array(27)(399),
      output(28) => mem_array(28)(399),
      output(29) => mem_array(29)(399),
      output(30) => mem_array(30)(399),
      output(31) => mem_array(31)(399),
      output(32) => mem_array(32)(399),
      output(33) => mem_array(33)(399),
      output(34) => mem_array(34)(399),
      output(35) => mem_array(35)(399)
      );
  rom400 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(400),
      output(0)  => mem_array(0)(400),
      output(1)  => mem_array(1)(400),
      output(2)  => mem_array(2)(400),
      output(3)  => mem_array(3)(400),
      output(4)  => mem_array(4)(400),
      output(5)  => mem_array(5)(400),
      output(6)  => mem_array(6)(400),
      output(7)  => mem_array(7)(400),
      output(8)  => mem_array(8)(400),
      output(9)  => mem_array(9)(400),
      output(10) => mem_array(10)(400),
      output(11) => mem_array(11)(400),
      output(12) => mem_array(12)(400),
      output(13) => mem_array(13)(400),
      output(14) => mem_array(14)(400),
      output(15) => mem_array(15)(400),
      output(16) => mem_array(16)(400),
      output(17) => mem_array(17)(400),
      output(18) => mem_array(18)(400),
      output(19) => mem_array(19)(400),
      output(20) => mem_array(20)(400),
      output(21) => mem_array(21)(400),
      output(22) => mem_array(22)(400),
      output(23) => mem_array(23)(400),
      output(24) => mem_array(24)(400),
      output(25) => mem_array(25)(400),
      output(26) => mem_array(26)(400),
      output(27) => mem_array(27)(400),
      output(28) => mem_array(28)(400),
      output(29) => mem_array(29)(400),
      output(30) => mem_array(30)(400),
      output(31) => mem_array(31)(400),
      output(32) => mem_array(32)(400),
      output(33) => mem_array(33)(400),
      output(34) => mem_array(34)(400),
      output(35) => mem_array(35)(400)
      );
  rom401 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(401),
      output(0)  => mem_array(0)(401),
      output(1)  => mem_array(1)(401),
      output(2)  => mem_array(2)(401),
      output(3)  => mem_array(3)(401),
      output(4)  => mem_array(4)(401),
      output(5)  => mem_array(5)(401),
      output(6)  => mem_array(6)(401),
      output(7)  => mem_array(7)(401),
      output(8)  => mem_array(8)(401),
      output(9)  => mem_array(9)(401),
      output(10) => mem_array(10)(401),
      output(11) => mem_array(11)(401),
      output(12) => mem_array(12)(401),
      output(13) => mem_array(13)(401),
      output(14) => mem_array(14)(401),
      output(15) => mem_array(15)(401),
      output(16) => mem_array(16)(401),
      output(17) => mem_array(17)(401),
      output(18) => mem_array(18)(401),
      output(19) => mem_array(19)(401),
      output(20) => mem_array(20)(401),
      output(21) => mem_array(21)(401),
      output(22) => mem_array(22)(401),
      output(23) => mem_array(23)(401),
      output(24) => mem_array(24)(401),
      output(25) => mem_array(25)(401),
      output(26) => mem_array(26)(401),
      output(27) => mem_array(27)(401),
      output(28) => mem_array(28)(401),
      output(29) => mem_array(29)(401),
      output(30) => mem_array(30)(401),
      output(31) => mem_array(31)(401),
      output(32) => mem_array(32)(401),
      output(33) => mem_array(33)(401),
      output(34) => mem_array(34)(401),
      output(35) => mem_array(35)(401)
      );
  rom402 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(402),
      output(0)  => mem_array(0)(402),
      output(1)  => mem_array(1)(402),
      output(2)  => mem_array(2)(402),
      output(3)  => mem_array(3)(402),
      output(4)  => mem_array(4)(402),
      output(5)  => mem_array(5)(402),
      output(6)  => mem_array(6)(402),
      output(7)  => mem_array(7)(402),
      output(8)  => mem_array(8)(402),
      output(9)  => mem_array(9)(402),
      output(10) => mem_array(10)(402),
      output(11) => mem_array(11)(402),
      output(12) => mem_array(12)(402),
      output(13) => mem_array(13)(402),
      output(14) => mem_array(14)(402),
      output(15) => mem_array(15)(402),
      output(16) => mem_array(16)(402),
      output(17) => mem_array(17)(402),
      output(18) => mem_array(18)(402),
      output(19) => mem_array(19)(402),
      output(20) => mem_array(20)(402),
      output(21) => mem_array(21)(402),
      output(22) => mem_array(22)(402),
      output(23) => mem_array(23)(402),
      output(24) => mem_array(24)(402),
      output(25) => mem_array(25)(402),
      output(26) => mem_array(26)(402),
      output(27) => mem_array(27)(402),
      output(28) => mem_array(28)(402),
      output(29) => mem_array(29)(402),
      output(30) => mem_array(30)(402),
      output(31) => mem_array(31)(402),
      output(32) => mem_array(32)(402),
      output(33) => mem_array(33)(402),
      output(34) => mem_array(34)(402),
      output(35) => mem_array(35)(402)
      );
  rom403 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(403),
      output(0)  => mem_array(0)(403),
      output(1)  => mem_array(1)(403),
      output(2)  => mem_array(2)(403),
      output(3)  => mem_array(3)(403),
      output(4)  => mem_array(4)(403),
      output(5)  => mem_array(5)(403),
      output(6)  => mem_array(6)(403),
      output(7)  => mem_array(7)(403),
      output(8)  => mem_array(8)(403),
      output(9)  => mem_array(9)(403),
      output(10) => mem_array(10)(403),
      output(11) => mem_array(11)(403),
      output(12) => mem_array(12)(403),
      output(13) => mem_array(13)(403),
      output(14) => mem_array(14)(403),
      output(15) => mem_array(15)(403),
      output(16) => mem_array(16)(403),
      output(17) => mem_array(17)(403),
      output(18) => mem_array(18)(403),
      output(19) => mem_array(19)(403),
      output(20) => mem_array(20)(403),
      output(21) => mem_array(21)(403),
      output(22) => mem_array(22)(403),
      output(23) => mem_array(23)(403),
      output(24) => mem_array(24)(403),
      output(25) => mem_array(25)(403),
      output(26) => mem_array(26)(403),
      output(27) => mem_array(27)(403),
      output(28) => mem_array(28)(403),
      output(29) => mem_array(29)(403),
      output(30) => mem_array(30)(403),
      output(31) => mem_array(31)(403),
      output(32) => mem_array(32)(403),
      output(33) => mem_array(33)(403),
      output(34) => mem_array(34)(403),
      output(35) => mem_array(35)(403)
      );
  rom404 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(404),
      output(0)  => mem_array(0)(404),
      output(1)  => mem_array(1)(404),
      output(2)  => mem_array(2)(404),
      output(3)  => mem_array(3)(404),
      output(4)  => mem_array(4)(404),
      output(5)  => mem_array(5)(404),
      output(6)  => mem_array(6)(404),
      output(7)  => mem_array(7)(404),
      output(8)  => mem_array(8)(404),
      output(9)  => mem_array(9)(404),
      output(10) => mem_array(10)(404),
      output(11) => mem_array(11)(404),
      output(12) => mem_array(12)(404),
      output(13) => mem_array(13)(404),
      output(14) => mem_array(14)(404),
      output(15) => mem_array(15)(404),
      output(16) => mem_array(16)(404),
      output(17) => mem_array(17)(404),
      output(18) => mem_array(18)(404),
      output(19) => mem_array(19)(404),
      output(20) => mem_array(20)(404),
      output(21) => mem_array(21)(404),
      output(22) => mem_array(22)(404),
      output(23) => mem_array(23)(404),
      output(24) => mem_array(24)(404),
      output(25) => mem_array(25)(404),
      output(26) => mem_array(26)(404),
      output(27) => mem_array(27)(404),
      output(28) => mem_array(28)(404),
      output(29) => mem_array(29)(404),
      output(30) => mem_array(30)(404),
      output(31) => mem_array(31)(404),
      output(32) => mem_array(32)(404),
      output(33) => mem_array(33)(404),
      output(34) => mem_array(34)(404),
      output(35) => mem_array(35)(404)
      );
  rom405 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(405),
      output(0)  => mem_array(0)(405),
      output(1)  => mem_array(1)(405),
      output(2)  => mem_array(2)(405),
      output(3)  => mem_array(3)(405),
      output(4)  => mem_array(4)(405),
      output(5)  => mem_array(5)(405),
      output(6)  => mem_array(6)(405),
      output(7)  => mem_array(7)(405),
      output(8)  => mem_array(8)(405),
      output(9)  => mem_array(9)(405),
      output(10) => mem_array(10)(405),
      output(11) => mem_array(11)(405),
      output(12) => mem_array(12)(405),
      output(13) => mem_array(13)(405),
      output(14) => mem_array(14)(405),
      output(15) => mem_array(15)(405),
      output(16) => mem_array(16)(405),
      output(17) => mem_array(17)(405),
      output(18) => mem_array(18)(405),
      output(19) => mem_array(19)(405),
      output(20) => mem_array(20)(405),
      output(21) => mem_array(21)(405),
      output(22) => mem_array(22)(405),
      output(23) => mem_array(23)(405),
      output(24) => mem_array(24)(405),
      output(25) => mem_array(25)(405),
      output(26) => mem_array(26)(405),
      output(27) => mem_array(27)(405),
      output(28) => mem_array(28)(405),
      output(29) => mem_array(29)(405),
      output(30) => mem_array(30)(405),
      output(31) => mem_array(31)(405),
      output(32) => mem_array(32)(405),
      output(33) => mem_array(33)(405),
      output(34) => mem_array(34)(405),
      output(35) => mem_array(35)(405)
      );
  rom406 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(406),
      output(0)  => mem_array(0)(406),
      output(1)  => mem_array(1)(406),
      output(2)  => mem_array(2)(406),
      output(3)  => mem_array(3)(406),
      output(4)  => mem_array(4)(406),
      output(5)  => mem_array(5)(406),
      output(6)  => mem_array(6)(406),
      output(7)  => mem_array(7)(406),
      output(8)  => mem_array(8)(406),
      output(9)  => mem_array(9)(406),
      output(10) => mem_array(10)(406),
      output(11) => mem_array(11)(406),
      output(12) => mem_array(12)(406),
      output(13) => mem_array(13)(406),
      output(14) => mem_array(14)(406),
      output(15) => mem_array(15)(406),
      output(16) => mem_array(16)(406),
      output(17) => mem_array(17)(406),
      output(18) => mem_array(18)(406),
      output(19) => mem_array(19)(406),
      output(20) => mem_array(20)(406),
      output(21) => mem_array(21)(406),
      output(22) => mem_array(22)(406),
      output(23) => mem_array(23)(406),
      output(24) => mem_array(24)(406),
      output(25) => mem_array(25)(406),
      output(26) => mem_array(26)(406),
      output(27) => mem_array(27)(406),
      output(28) => mem_array(28)(406),
      output(29) => mem_array(29)(406),
      output(30) => mem_array(30)(406),
      output(31) => mem_array(31)(406),
      output(32) => mem_array(32)(406),
      output(33) => mem_array(33)(406),
      output(34) => mem_array(34)(406),
      output(35) => mem_array(35)(406)
      );
  rom407 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(407),
      output(0)  => mem_array(0)(407),
      output(1)  => mem_array(1)(407),
      output(2)  => mem_array(2)(407),
      output(3)  => mem_array(3)(407),
      output(4)  => mem_array(4)(407),
      output(5)  => mem_array(5)(407),
      output(6)  => mem_array(6)(407),
      output(7)  => mem_array(7)(407),
      output(8)  => mem_array(8)(407),
      output(9)  => mem_array(9)(407),
      output(10) => mem_array(10)(407),
      output(11) => mem_array(11)(407),
      output(12) => mem_array(12)(407),
      output(13) => mem_array(13)(407),
      output(14) => mem_array(14)(407),
      output(15) => mem_array(15)(407),
      output(16) => mem_array(16)(407),
      output(17) => mem_array(17)(407),
      output(18) => mem_array(18)(407),
      output(19) => mem_array(19)(407),
      output(20) => mem_array(20)(407),
      output(21) => mem_array(21)(407),
      output(22) => mem_array(22)(407),
      output(23) => mem_array(23)(407),
      output(24) => mem_array(24)(407),
      output(25) => mem_array(25)(407),
      output(26) => mem_array(26)(407),
      output(27) => mem_array(27)(407),
      output(28) => mem_array(28)(407),
      output(29) => mem_array(29)(407),
      output(30) => mem_array(30)(407),
      output(31) => mem_array(31)(407),
      output(32) => mem_array(32)(407),
      output(33) => mem_array(33)(407),
      output(34) => mem_array(34)(407),
      output(35) => mem_array(35)(407)
      );
  rom408 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(408),
      output(0)  => mem_array(0)(408),
      output(1)  => mem_array(1)(408),
      output(2)  => mem_array(2)(408),
      output(3)  => mem_array(3)(408),
      output(4)  => mem_array(4)(408),
      output(5)  => mem_array(5)(408),
      output(6)  => mem_array(6)(408),
      output(7)  => mem_array(7)(408),
      output(8)  => mem_array(8)(408),
      output(9)  => mem_array(9)(408),
      output(10) => mem_array(10)(408),
      output(11) => mem_array(11)(408),
      output(12) => mem_array(12)(408),
      output(13) => mem_array(13)(408),
      output(14) => mem_array(14)(408),
      output(15) => mem_array(15)(408),
      output(16) => mem_array(16)(408),
      output(17) => mem_array(17)(408),
      output(18) => mem_array(18)(408),
      output(19) => mem_array(19)(408),
      output(20) => mem_array(20)(408),
      output(21) => mem_array(21)(408),
      output(22) => mem_array(22)(408),
      output(23) => mem_array(23)(408),
      output(24) => mem_array(24)(408),
      output(25) => mem_array(25)(408),
      output(26) => mem_array(26)(408),
      output(27) => mem_array(27)(408),
      output(28) => mem_array(28)(408),
      output(29) => mem_array(29)(408),
      output(30) => mem_array(30)(408),
      output(31) => mem_array(31)(408),
      output(32) => mem_array(32)(408),
      output(33) => mem_array(33)(408),
      output(34) => mem_array(34)(408),
      output(35) => mem_array(35)(408)
      );
  rom409 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(409),
      output(0)  => mem_array(0)(409),
      output(1)  => mem_array(1)(409),
      output(2)  => mem_array(2)(409),
      output(3)  => mem_array(3)(409),
      output(4)  => mem_array(4)(409),
      output(5)  => mem_array(5)(409),
      output(6)  => mem_array(6)(409),
      output(7)  => mem_array(7)(409),
      output(8)  => mem_array(8)(409),
      output(9)  => mem_array(9)(409),
      output(10) => mem_array(10)(409),
      output(11) => mem_array(11)(409),
      output(12) => mem_array(12)(409),
      output(13) => mem_array(13)(409),
      output(14) => mem_array(14)(409),
      output(15) => mem_array(15)(409),
      output(16) => mem_array(16)(409),
      output(17) => mem_array(17)(409),
      output(18) => mem_array(18)(409),
      output(19) => mem_array(19)(409),
      output(20) => mem_array(20)(409),
      output(21) => mem_array(21)(409),
      output(22) => mem_array(22)(409),
      output(23) => mem_array(23)(409),
      output(24) => mem_array(24)(409),
      output(25) => mem_array(25)(409),
      output(26) => mem_array(26)(409),
      output(27) => mem_array(27)(409),
      output(28) => mem_array(28)(409),
      output(29) => mem_array(29)(409),
      output(30) => mem_array(30)(409),
      output(31) => mem_array(31)(409),
      output(32) => mem_array(32)(409),
      output(33) => mem_array(33)(409),
      output(34) => mem_array(34)(409),
      output(35) => mem_array(35)(409)
      );
  rom410 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(410),
      output(0)  => mem_array(0)(410),
      output(1)  => mem_array(1)(410),
      output(2)  => mem_array(2)(410),
      output(3)  => mem_array(3)(410),
      output(4)  => mem_array(4)(410),
      output(5)  => mem_array(5)(410),
      output(6)  => mem_array(6)(410),
      output(7)  => mem_array(7)(410),
      output(8)  => mem_array(8)(410),
      output(9)  => mem_array(9)(410),
      output(10) => mem_array(10)(410),
      output(11) => mem_array(11)(410),
      output(12) => mem_array(12)(410),
      output(13) => mem_array(13)(410),
      output(14) => mem_array(14)(410),
      output(15) => mem_array(15)(410),
      output(16) => mem_array(16)(410),
      output(17) => mem_array(17)(410),
      output(18) => mem_array(18)(410),
      output(19) => mem_array(19)(410),
      output(20) => mem_array(20)(410),
      output(21) => mem_array(21)(410),
      output(22) => mem_array(22)(410),
      output(23) => mem_array(23)(410),
      output(24) => mem_array(24)(410),
      output(25) => mem_array(25)(410),
      output(26) => mem_array(26)(410),
      output(27) => mem_array(27)(410),
      output(28) => mem_array(28)(410),
      output(29) => mem_array(29)(410),
      output(30) => mem_array(30)(410),
      output(31) => mem_array(31)(410),
      output(32) => mem_array(32)(410),
      output(33) => mem_array(33)(410),
      output(34) => mem_array(34)(410),
      output(35) => mem_array(35)(410)
      );
  rom411 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(411),
      output(0)  => mem_array(0)(411),
      output(1)  => mem_array(1)(411),
      output(2)  => mem_array(2)(411),
      output(3)  => mem_array(3)(411),
      output(4)  => mem_array(4)(411),
      output(5)  => mem_array(5)(411),
      output(6)  => mem_array(6)(411),
      output(7)  => mem_array(7)(411),
      output(8)  => mem_array(8)(411),
      output(9)  => mem_array(9)(411),
      output(10) => mem_array(10)(411),
      output(11) => mem_array(11)(411),
      output(12) => mem_array(12)(411),
      output(13) => mem_array(13)(411),
      output(14) => mem_array(14)(411),
      output(15) => mem_array(15)(411),
      output(16) => mem_array(16)(411),
      output(17) => mem_array(17)(411),
      output(18) => mem_array(18)(411),
      output(19) => mem_array(19)(411),
      output(20) => mem_array(20)(411),
      output(21) => mem_array(21)(411),
      output(22) => mem_array(22)(411),
      output(23) => mem_array(23)(411),
      output(24) => mem_array(24)(411),
      output(25) => mem_array(25)(411),
      output(26) => mem_array(26)(411),
      output(27) => mem_array(27)(411),
      output(28) => mem_array(28)(411),
      output(29) => mem_array(29)(411),
      output(30) => mem_array(30)(411),
      output(31) => mem_array(31)(411),
      output(32) => mem_array(32)(411),
      output(33) => mem_array(33)(411),
      output(34) => mem_array(34)(411),
      output(35) => mem_array(35)(411)
      );
  rom412 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(412),
      output(0)  => mem_array(0)(412),
      output(1)  => mem_array(1)(412),
      output(2)  => mem_array(2)(412),
      output(3)  => mem_array(3)(412),
      output(4)  => mem_array(4)(412),
      output(5)  => mem_array(5)(412),
      output(6)  => mem_array(6)(412),
      output(7)  => mem_array(7)(412),
      output(8)  => mem_array(8)(412),
      output(9)  => mem_array(9)(412),
      output(10) => mem_array(10)(412),
      output(11) => mem_array(11)(412),
      output(12) => mem_array(12)(412),
      output(13) => mem_array(13)(412),
      output(14) => mem_array(14)(412),
      output(15) => mem_array(15)(412),
      output(16) => mem_array(16)(412),
      output(17) => mem_array(17)(412),
      output(18) => mem_array(18)(412),
      output(19) => mem_array(19)(412),
      output(20) => mem_array(20)(412),
      output(21) => mem_array(21)(412),
      output(22) => mem_array(22)(412),
      output(23) => mem_array(23)(412),
      output(24) => mem_array(24)(412),
      output(25) => mem_array(25)(412),
      output(26) => mem_array(26)(412),
      output(27) => mem_array(27)(412),
      output(28) => mem_array(28)(412),
      output(29) => mem_array(29)(412),
      output(30) => mem_array(30)(412),
      output(31) => mem_array(31)(412),
      output(32) => mem_array(32)(412),
      output(33) => mem_array(33)(412),
      output(34) => mem_array(34)(412),
      output(35) => mem_array(35)(412)
      );
  rom413 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(413),
      output(0)  => mem_array(0)(413),
      output(1)  => mem_array(1)(413),
      output(2)  => mem_array(2)(413),
      output(3)  => mem_array(3)(413),
      output(4)  => mem_array(4)(413),
      output(5)  => mem_array(5)(413),
      output(6)  => mem_array(6)(413),
      output(7)  => mem_array(7)(413),
      output(8)  => mem_array(8)(413),
      output(9)  => mem_array(9)(413),
      output(10) => mem_array(10)(413),
      output(11) => mem_array(11)(413),
      output(12) => mem_array(12)(413),
      output(13) => mem_array(13)(413),
      output(14) => mem_array(14)(413),
      output(15) => mem_array(15)(413),
      output(16) => mem_array(16)(413),
      output(17) => mem_array(17)(413),
      output(18) => mem_array(18)(413),
      output(19) => mem_array(19)(413),
      output(20) => mem_array(20)(413),
      output(21) => mem_array(21)(413),
      output(22) => mem_array(22)(413),
      output(23) => mem_array(23)(413),
      output(24) => mem_array(24)(413),
      output(25) => mem_array(25)(413),
      output(26) => mem_array(26)(413),
      output(27) => mem_array(27)(413),
      output(28) => mem_array(28)(413),
      output(29) => mem_array(29)(413),
      output(30) => mem_array(30)(413),
      output(31) => mem_array(31)(413),
      output(32) => mem_array(32)(413),
      output(33) => mem_array(33)(413),
      output(34) => mem_array(34)(413),
      output(35) => mem_array(35)(413)
      );
  rom414 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(414),
      output(0)  => mem_array(0)(414),
      output(1)  => mem_array(1)(414),
      output(2)  => mem_array(2)(414),
      output(3)  => mem_array(3)(414),
      output(4)  => mem_array(4)(414),
      output(5)  => mem_array(5)(414),
      output(6)  => mem_array(6)(414),
      output(7)  => mem_array(7)(414),
      output(8)  => mem_array(8)(414),
      output(9)  => mem_array(9)(414),
      output(10) => mem_array(10)(414),
      output(11) => mem_array(11)(414),
      output(12) => mem_array(12)(414),
      output(13) => mem_array(13)(414),
      output(14) => mem_array(14)(414),
      output(15) => mem_array(15)(414),
      output(16) => mem_array(16)(414),
      output(17) => mem_array(17)(414),
      output(18) => mem_array(18)(414),
      output(19) => mem_array(19)(414),
      output(20) => mem_array(20)(414),
      output(21) => mem_array(21)(414),
      output(22) => mem_array(22)(414),
      output(23) => mem_array(23)(414),
      output(24) => mem_array(24)(414),
      output(25) => mem_array(25)(414),
      output(26) => mem_array(26)(414),
      output(27) => mem_array(27)(414),
      output(28) => mem_array(28)(414),
      output(29) => mem_array(29)(414),
      output(30) => mem_array(30)(414),
      output(31) => mem_array(31)(414),
      output(32) => mem_array(32)(414),
      output(33) => mem_array(33)(414),
      output(34) => mem_array(34)(414),
      output(35) => mem_array(35)(414)
      );
  rom415 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(415),
      output(0)  => mem_array(0)(415),
      output(1)  => mem_array(1)(415),
      output(2)  => mem_array(2)(415),
      output(3)  => mem_array(3)(415),
      output(4)  => mem_array(4)(415),
      output(5)  => mem_array(5)(415),
      output(6)  => mem_array(6)(415),
      output(7)  => mem_array(7)(415),
      output(8)  => mem_array(8)(415),
      output(9)  => mem_array(9)(415),
      output(10) => mem_array(10)(415),
      output(11) => mem_array(11)(415),
      output(12) => mem_array(12)(415),
      output(13) => mem_array(13)(415),
      output(14) => mem_array(14)(415),
      output(15) => mem_array(15)(415),
      output(16) => mem_array(16)(415),
      output(17) => mem_array(17)(415),
      output(18) => mem_array(18)(415),
      output(19) => mem_array(19)(415),
      output(20) => mem_array(20)(415),
      output(21) => mem_array(21)(415),
      output(22) => mem_array(22)(415),
      output(23) => mem_array(23)(415),
      output(24) => mem_array(24)(415),
      output(25) => mem_array(25)(415),
      output(26) => mem_array(26)(415),
      output(27) => mem_array(27)(415),
      output(28) => mem_array(28)(415),
      output(29) => mem_array(29)(415),
      output(30) => mem_array(30)(415),
      output(31) => mem_array(31)(415),
      output(32) => mem_array(32)(415),
      output(33) => mem_array(33)(415),
      output(34) => mem_array(34)(415),
      output(35) => mem_array(35)(415)
      );
  rom416 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(416),
      output(0)  => mem_array(0)(416),
      output(1)  => mem_array(1)(416),
      output(2)  => mem_array(2)(416),
      output(3)  => mem_array(3)(416),
      output(4)  => mem_array(4)(416),
      output(5)  => mem_array(5)(416),
      output(6)  => mem_array(6)(416),
      output(7)  => mem_array(7)(416),
      output(8)  => mem_array(8)(416),
      output(9)  => mem_array(9)(416),
      output(10) => mem_array(10)(416),
      output(11) => mem_array(11)(416),
      output(12) => mem_array(12)(416),
      output(13) => mem_array(13)(416),
      output(14) => mem_array(14)(416),
      output(15) => mem_array(15)(416),
      output(16) => mem_array(16)(416),
      output(17) => mem_array(17)(416),
      output(18) => mem_array(18)(416),
      output(19) => mem_array(19)(416),
      output(20) => mem_array(20)(416),
      output(21) => mem_array(21)(416),
      output(22) => mem_array(22)(416),
      output(23) => mem_array(23)(416),
      output(24) => mem_array(24)(416),
      output(25) => mem_array(25)(416),
      output(26) => mem_array(26)(416),
      output(27) => mem_array(27)(416),
      output(28) => mem_array(28)(416),
      output(29) => mem_array(29)(416),
      output(30) => mem_array(30)(416),
      output(31) => mem_array(31)(416),
      output(32) => mem_array(32)(416),
      output(33) => mem_array(33)(416),
      output(34) => mem_array(34)(416),
      output(35) => mem_array(35)(416)
      );
  rom417 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(417),
      output(0)  => mem_array(0)(417),
      output(1)  => mem_array(1)(417),
      output(2)  => mem_array(2)(417),
      output(3)  => mem_array(3)(417),
      output(4)  => mem_array(4)(417),
      output(5)  => mem_array(5)(417),
      output(6)  => mem_array(6)(417),
      output(7)  => mem_array(7)(417),
      output(8)  => mem_array(8)(417),
      output(9)  => mem_array(9)(417),
      output(10) => mem_array(10)(417),
      output(11) => mem_array(11)(417),
      output(12) => mem_array(12)(417),
      output(13) => mem_array(13)(417),
      output(14) => mem_array(14)(417),
      output(15) => mem_array(15)(417),
      output(16) => mem_array(16)(417),
      output(17) => mem_array(17)(417),
      output(18) => mem_array(18)(417),
      output(19) => mem_array(19)(417),
      output(20) => mem_array(20)(417),
      output(21) => mem_array(21)(417),
      output(22) => mem_array(22)(417),
      output(23) => mem_array(23)(417),
      output(24) => mem_array(24)(417),
      output(25) => mem_array(25)(417),
      output(26) => mem_array(26)(417),
      output(27) => mem_array(27)(417),
      output(28) => mem_array(28)(417),
      output(29) => mem_array(29)(417),
      output(30) => mem_array(30)(417),
      output(31) => mem_array(31)(417),
      output(32) => mem_array(32)(417),
      output(33) => mem_array(33)(417),
      output(34) => mem_array(34)(417),
      output(35) => mem_array(35)(417)
      );
  rom418 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(418),
      output(0)  => mem_array(0)(418),
      output(1)  => mem_array(1)(418),
      output(2)  => mem_array(2)(418),
      output(3)  => mem_array(3)(418),
      output(4)  => mem_array(4)(418),
      output(5)  => mem_array(5)(418),
      output(6)  => mem_array(6)(418),
      output(7)  => mem_array(7)(418),
      output(8)  => mem_array(8)(418),
      output(9)  => mem_array(9)(418),
      output(10) => mem_array(10)(418),
      output(11) => mem_array(11)(418),
      output(12) => mem_array(12)(418),
      output(13) => mem_array(13)(418),
      output(14) => mem_array(14)(418),
      output(15) => mem_array(15)(418),
      output(16) => mem_array(16)(418),
      output(17) => mem_array(17)(418),
      output(18) => mem_array(18)(418),
      output(19) => mem_array(19)(418),
      output(20) => mem_array(20)(418),
      output(21) => mem_array(21)(418),
      output(22) => mem_array(22)(418),
      output(23) => mem_array(23)(418),
      output(24) => mem_array(24)(418),
      output(25) => mem_array(25)(418),
      output(26) => mem_array(26)(418),
      output(27) => mem_array(27)(418),
      output(28) => mem_array(28)(418),
      output(29) => mem_array(29)(418),
      output(30) => mem_array(30)(418),
      output(31) => mem_array(31)(418),
      output(32) => mem_array(32)(418),
      output(33) => mem_array(33)(418),
      output(34) => mem_array(34)(418),
      output(35) => mem_array(35)(418)
      );
  rom419 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(419),
      output(0)  => mem_array(0)(419),
      output(1)  => mem_array(1)(419),
      output(2)  => mem_array(2)(419),
      output(3)  => mem_array(3)(419),
      output(4)  => mem_array(4)(419),
      output(5)  => mem_array(5)(419),
      output(6)  => mem_array(6)(419),
      output(7)  => mem_array(7)(419),
      output(8)  => mem_array(8)(419),
      output(9)  => mem_array(9)(419),
      output(10) => mem_array(10)(419),
      output(11) => mem_array(11)(419),
      output(12) => mem_array(12)(419),
      output(13) => mem_array(13)(419),
      output(14) => mem_array(14)(419),
      output(15) => mem_array(15)(419),
      output(16) => mem_array(16)(419),
      output(17) => mem_array(17)(419),
      output(18) => mem_array(18)(419),
      output(19) => mem_array(19)(419),
      output(20) => mem_array(20)(419),
      output(21) => mem_array(21)(419),
      output(22) => mem_array(22)(419),
      output(23) => mem_array(23)(419),
      output(24) => mem_array(24)(419),
      output(25) => mem_array(25)(419),
      output(26) => mem_array(26)(419),
      output(27) => mem_array(27)(419),
      output(28) => mem_array(28)(419),
      output(29) => mem_array(29)(419),
      output(30) => mem_array(30)(419),
      output(31) => mem_array(31)(419),
      output(32) => mem_array(32)(419),
      output(33) => mem_array(33)(419),
      output(34) => mem_array(34)(419),
      output(35) => mem_array(35)(419)
      );
  rom420 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(420),
      output(0)  => mem_array(0)(420),
      output(1)  => mem_array(1)(420),
      output(2)  => mem_array(2)(420),
      output(3)  => mem_array(3)(420),
      output(4)  => mem_array(4)(420),
      output(5)  => mem_array(5)(420),
      output(6)  => mem_array(6)(420),
      output(7)  => mem_array(7)(420),
      output(8)  => mem_array(8)(420),
      output(9)  => mem_array(9)(420),
      output(10) => mem_array(10)(420),
      output(11) => mem_array(11)(420),
      output(12) => mem_array(12)(420),
      output(13) => mem_array(13)(420),
      output(14) => mem_array(14)(420),
      output(15) => mem_array(15)(420),
      output(16) => mem_array(16)(420),
      output(17) => mem_array(17)(420),
      output(18) => mem_array(18)(420),
      output(19) => mem_array(19)(420),
      output(20) => mem_array(20)(420),
      output(21) => mem_array(21)(420),
      output(22) => mem_array(22)(420),
      output(23) => mem_array(23)(420),
      output(24) => mem_array(24)(420),
      output(25) => mem_array(25)(420),
      output(26) => mem_array(26)(420),
      output(27) => mem_array(27)(420),
      output(28) => mem_array(28)(420),
      output(29) => mem_array(29)(420),
      output(30) => mem_array(30)(420),
      output(31) => mem_array(31)(420),
      output(32) => mem_array(32)(420),
      output(33) => mem_array(33)(420),
      output(34) => mem_array(34)(420),
      output(35) => mem_array(35)(420)
      );
  rom421 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(421),
      output(0)  => mem_array(0)(421),
      output(1)  => mem_array(1)(421),
      output(2)  => mem_array(2)(421),
      output(3)  => mem_array(3)(421),
      output(4)  => mem_array(4)(421),
      output(5)  => mem_array(5)(421),
      output(6)  => mem_array(6)(421),
      output(7)  => mem_array(7)(421),
      output(8)  => mem_array(8)(421),
      output(9)  => mem_array(9)(421),
      output(10) => mem_array(10)(421),
      output(11) => mem_array(11)(421),
      output(12) => mem_array(12)(421),
      output(13) => mem_array(13)(421),
      output(14) => mem_array(14)(421),
      output(15) => mem_array(15)(421),
      output(16) => mem_array(16)(421),
      output(17) => mem_array(17)(421),
      output(18) => mem_array(18)(421),
      output(19) => mem_array(19)(421),
      output(20) => mem_array(20)(421),
      output(21) => mem_array(21)(421),
      output(22) => mem_array(22)(421),
      output(23) => mem_array(23)(421),
      output(24) => mem_array(24)(421),
      output(25) => mem_array(25)(421),
      output(26) => mem_array(26)(421),
      output(27) => mem_array(27)(421),
      output(28) => mem_array(28)(421),
      output(29) => mem_array(29)(421),
      output(30) => mem_array(30)(421),
      output(31) => mem_array(31)(421),
      output(32) => mem_array(32)(421),
      output(33) => mem_array(33)(421),
      output(34) => mem_array(34)(421),
      output(35) => mem_array(35)(421)
      );
  rom422 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(422),
      output(0)  => mem_array(0)(422),
      output(1)  => mem_array(1)(422),
      output(2)  => mem_array(2)(422),
      output(3)  => mem_array(3)(422),
      output(4)  => mem_array(4)(422),
      output(5)  => mem_array(5)(422),
      output(6)  => mem_array(6)(422),
      output(7)  => mem_array(7)(422),
      output(8)  => mem_array(8)(422),
      output(9)  => mem_array(9)(422),
      output(10) => mem_array(10)(422),
      output(11) => mem_array(11)(422),
      output(12) => mem_array(12)(422),
      output(13) => mem_array(13)(422),
      output(14) => mem_array(14)(422),
      output(15) => mem_array(15)(422),
      output(16) => mem_array(16)(422),
      output(17) => mem_array(17)(422),
      output(18) => mem_array(18)(422),
      output(19) => mem_array(19)(422),
      output(20) => mem_array(20)(422),
      output(21) => mem_array(21)(422),
      output(22) => mem_array(22)(422),
      output(23) => mem_array(23)(422),
      output(24) => mem_array(24)(422),
      output(25) => mem_array(25)(422),
      output(26) => mem_array(26)(422),
      output(27) => mem_array(27)(422),
      output(28) => mem_array(28)(422),
      output(29) => mem_array(29)(422),
      output(30) => mem_array(30)(422),
      output(31) => mem_array(31)(422),
      output(32) => mem_array(32)(422),
      output(33) => mem_array(33)(422),
      output(34) => mem_array(34)(422),
      output(35) => mem_array(35)(422)
      );
  rom423 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(423),
      output(0)  => mem_array(0)(423),
      output(1)  => mem_array(1)(423),
      output(2)  => mem_array(2)(423),
      output(3)  => mem_array(3)(423),
      output(4)  => mem_array(4)(423),
      output(5)  => mem_array(5)(423),
      output(6)  => mem_array(6)(423),
      output(7)  => mem_array(7)(423),
      output(8)  => mem_array(8)(423),
      output(9)  => mem_array(9)(423),
      output(10) => mem_array(10)(423),
      output(11) => mem_array(11)(423),
      output(12) => mem_array(12)(423),
      output(13) => mem_array(13)(423),
      output(14) => mem_array(14)(423),
      output(15) => mem_array(15)(423),
      output(16) => mem_array(16)(423),
      output(17) => mem_array(17)(423),
      output(18) => mem_array(18)(423),
      output(19) => mem_array(19)(423),
      output(20) => mem_array(20)(423),
      output(21) => mem_array(21)(423),
      output(22) => mem_array(22)(423),
      output(23) => mem_array(23)(423),
      output(24) => mem_array(24)(423),
      output(25) => mem_array(25)(423),
      output(26) => mem_array(26)(423),
      output(27) => mem_array(27)(423),
      output(28) => mem_array(28)(423),
      output(29) => mem_array(29)(423),
      output(30) => mem_array(30)(423),
      output(31) => mem_array(31)(423),
      output(32) => mem_array(32)(423),
      output(33) => mem_array(33)(423),
      output(34) => mem_array(34)(423),
      output(35) => mem_array(35)(423)
      );
  rom424 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(424),
      output(0)  => mem_array(0)(424),
      output(1)  => mem_array(1)(424),
      output(2)  => mem_array(2)(424),
      output(3)  => mem_array(3)(424),
      output(4)  => mem_array(4)(424),
      output(5)  => mem_array(5)(424),
      output(6)  => mem_array(6)(424),
      output(7)  => mem_array(7)(424),
      output(8)  => mem_array(8)(424),
      output(9)  => mem_array(9)(424),
      output(10) => mem_array(10)(424),
      output(11) => mem_array(11)(424),
      output(12) => mem_array(12)(424),
      output(13) => mem_array(13)(424),
      output(14) => mem_array(14)(424),
      output(15) => mem_array(15)(424),
      output(16) => mem_array(16)(424),
      output(17) => mem_array(17)(424),
      output(18) => mem_array(18)(424),
      output(19) => mem_array(19)(424),
      output(20) => mem_array(20)(424),
      output(21) => mem_array(21)(424),
      output(22) => mem_array(22)(424),
      output(23) => mem_array(23)(424),
      output(24) => mem_array(24)(424),
      output(25) => mem_array(25)(424),
      output(26) => mem_array(26)(424),
      output(27) => mem_array(27)(424),
      output(28) => mem_array(28)(424),
      output(29) => mem_array(29)(424),
      output(30) => mem_array(30)(424),
      output(31) => mem_array(31)(424),
      output(32) => mem_array(32)(424),
      output(33) => mem_array(33)(424),
      output(34) => mem_array(34)(424),
      output(35) => mem_array(35)(424)
      );
  rom425 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(425),
      output(0)  => mem_array(0)(425),
      output(1)  => mem_array(1)(425),
      output(2)  => mem_array(2)(425),
      output(3)  => mem_array(3)(425),
      output(4)  => mem_array(4)(425),
      output(5)  => mem_array(5)(425),
      output(6)  => mem_array(6)(425),
      output(7)  => mem_array(7)(425),
      output(8)  => mem_array(8)(425),
      output(9)  => mem_array(9)(425),
      output(10) => mem_array(10)(425),
      output(11) => mem_array(11)(425),
      output(12) => mem_array(12)(425),
      output(13) => mem_array(13)(425),
      output(14) => mem_array(14)(425),
      output(15) => mem_array(15)(425),
      output(16) => mem_array(16)(425),
      output(17) => mem_array(17)(425),
      output(18) => mem_array(18)(425),
      output(19) => mem_array(19)(425),
      output(20) => mem_array(20)(425),
      output(21) => mem_array(21)(425),
      output(22) => mem_array(22)(425),
      output(23) => mem_array(23)(425),
      output(24) => mem_array(24)(425),
      output(25) => mem_array(25)(425),
      output(26) => mem_array(26)(425),
      output(27) => mem_array(27)(425),
      output(28) => mem_array(28)(425),
      output(29) => mem_array(29)(425),
      output(30) => mem_array(30)(425),
      output(31) => mem_array(31)(425),
      output(32) => mem_array(32)(425),
      output(33) => mem_array(33)(425),
      output(34) => mem_array(34)(425),
      output(35) => mem_array(35)(425)
      );
  rom426 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(426),
      output(0)  => mem_array(0)(426),
      output(1)  => mem_array(1)(426),
      output(2)  => mem_array(2)(426),
      output(3)  => mem_array(3)(426),
      output(4)  => mem_array(4)(426),
      output(5)  => mem_array(5)(426),
      output(6)  => mem_array(6)(426),
      output(7)  => mem_array(7)(426),
      output(8)  => mem_array(8)(426),
      output(9)  => mem_array(9)(426),
      output(10) => mem_array(10)(426),
      output(11) => mem_array(11)(426),
      output(12) => mem_array(12)(426),
      output(13) => mem_array(13)(426),
      output(14) => mem_array(14)(426),
      output(15) => mem_array(15)(426),
      output(16) => mem_array(16)(426),
      output(17) => mem_array(17)(426),
      output(18) => mem_array(18)(426),
      output(19) => mem_array(19)(426),
      output(20) => mem_array(20)(426),
      output(21) => mem_array(21)(426),
      output(22) => mem_array(22)(426),
      output(23) => mem_array(23)(426),
      output(24) => mem_array(24)(426),
      output(25) => mem_array(25)(426),
      output(26) => mem_array(26)(426),
      output(27) => mem_array(27)(426),
      output(28) => mem_array(28)(426),
      output(29) => mem_array(29)(426),
      output(30) => mem_array(30)(426),
      output(31) => mem_array(31)(426),
      output(32) => mem_array(32)(426),
      output(33) => mem_array(33)(426),
      output(34) => mem_array(34)(426),
      output(35) => mem_array(35)(426)
      );
  rom427 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(427),
      output(0)  => mem_array(0)(427),
      output(1)  => mem_array(1)(427),
      output(2)  => mem_array(2)(427),
      output(3)  => mem_array(3)(427),
      output(4)  => mem_array(4)(427),
      output(5)  => mem_array(5)(427),
      output(6)  => mem_array(6)(427),
      output(7)  => mem_array(7)(427),
      output(8)  => mem_array(8)(427),
      output(9)  => mem_array(9)(427),
      output(10) => mem_array(10)(427),
      output(11) => mem_array(11)(427),
      output(12) => mem_array(12)(427),
      output(13) => mem_array(13)(427),
      output(14) => mem_array(14)(427),
      output(15) => mem_array(15)(427),
      output(16) => mem_array(16)(427),
      output(17) => mem_array(17)(427),
      output(18) => mem_array(18)(427),
      output(19) => mem_array(19)(427),
      output(20) => mem_array(20)(427),
      output(21) => mem_array(21)(427),
      output(22) => mem_array(22)(427),
      output(23) => mem_array(23)(427),
      output(24) => mem_array(24)(427),
      output(25) => mem_array(25)(427),
      output(26) => mem_array(26)(427),
      output(27) => mem_array(27)(427),
      output(28) => mem_array(28)(427),
      output(29) => mem_array(29)(427),
      output(30) => mem_array(30)(427),
      output(31) => mem_array(31)(427),
      output(32) => mem_array(32)(427),
      output(33) => mem_array(33)(427),
      output(34) => mem_array(34)(427),
      output(35) => mem_array(35)(427)
      );
  rom428 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(428),
      output(0)  => mem_array(0)(428),
      output(1)  => mem_array(1)(428),
      output(2)  => mem_array(2)(428),
      output(3)  => mem_array(3)(428),
      output(4)  => mem_array(4)(428),
      output(5)  => mem_array(5)(428),
      output(6)  => mem_array(6)(428),
      output(7)  => mem_array(7)(428),
      output(8)  => mem_array(8)(428),
      output(9)  => mem_array(9)(428),
      output(10) => mem_array(10)(428),
      output(11) => mem_array(11)(428),
      output(12) => mem_array(12)(428),
      output(13) => mem_array(13)(428),
      output(14) => mem_array(14)(428),
      output(15) => mem_array(15)(428),
      output(16) => mem_array(16)(428),
      output(17) => mem_array(17)(428),
      output(18) => mem_array(18)(428),
      output(19) => mem_array(19)(428),
      output(20) => mem_array(20)(428),
      output(21) => mem_array(21)(428),
      output(22) => mem_array(22)(428),
      output(23) => mem_array(23)(428),
      output(24) => mem_array(24)(428),
      output(25) => mem_array(25)(428),
      output(26) => mem_array(26)(428),
      output(27) => mem_array(27)(428),
      output(28) => mem_array(28)(428),
      output(29) => mem_array(29)(428),
      output(30) => mem_array(30)(428),
      output(31) => mem_array(31)(428),
      output(32) => mem_array(32)(428),
      output(33) => mem_array(33)(428),
      output(34) => mem_array(34)(428),
      output(35) => mem_array(35)(428)
      );
  rom429 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(429),
      output(0)  => mem_array(0)(429),
      output(1)  => mem_array(1)(429),
      output(2)  => mem_array(2)(429),
      output(3)  => mem_array(3)(429),
      output(4)  => mem_array(4)(429),
      output(5)  => mem_array(5)(429),
      output(6)  => mem_array(6)(429),
      output(7)  => mem_array(7)(429),
      output(8)  => mem_array(8)(429),
      output(9)  => mem_array(9)(429),
      output(10) => mem_array(10)(429),
      output(11) => mem_array(11)(429),
      output(12) => mem_array(12)(429),
      output(13) => mem_array(13)(429),
      output(14) => mem_array(14)(429),
      output(15) => mem_array(15)(429),
      output(16) => mem_array(16)(429),
      output(17) => mem_array(17)(429),
      output(18) => mem_array(18)(429),
      output(19) => mem_array(19)(429),
      output(20) => mem_array(20)(429),
      output(21) => mem_array(21)(429),
      output(22) => mem_array(22)(429),
      output(23) => mem_array(23)(429),
      output(24) => mem_array(24)(429),
      output(25) => mem_array(25)(429),
      output(26) => mem_array(26)(429),
      output(27) => mem_array(27)(429),
      output(28) => mem_array(28)(429),
      output(29) => mem_array(29)(429),
      output(30) => mem_array(30)(429),
      output(31) => mem_array(31)(429),
      output(32) => mem_array(32)(429),
      output(33) => mem_array(33)(429),
      output(34) => mem_array(34)(429),
      output(35) => mem_array(35)(429)
      );
  rom430 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(430),
      output(0)  => mem_array(0)(430),
      output(1)  => mem_array(1)(430),
      output(2)  => mem_array(2)(430),
      output(3)  => mem_array(3)(430),
      output(4)  => mem_array(4)(430),
      output(5)  => mem_array(5)(430),
      output(6)  => mem_array(6)(430),
      output(7)  => mem_array(7)(430),
      output(8)  => mem_array(8)(430),
      output(9)  => mem_array(9)(430),
      output(10) => mem_array(10)(430),
      output(11) => mem_array(11)(430),
      output(12) => mem_array(12)(430),
      output(13) => mem_array(13)(430),
      output(14) => mem_array(14)(430),
      output(15) => mem_array(15)(430),
      output(16) => mem_array(16)(430),
      output(17) => mem_array(17)(430),
      output(18) => mem_array(18)(430),
      output(19) => mem_array(19)(430),
      output(20) => mem_array(20)(430),
      output(21) => mem_array(21)(430),
      output(22) => mem_array(22)(430),
      output(23) => mem_array(23)(430),
      output(24) => mem_array(24)(430),
      output(25) => mem_array(25)(430),
      output(26) => mem_array(26)(430),
      output(27) => mem_array(27)(430),
      output(28) => mem_array(28)(430),
      output(29) => mem_array(29)(430),
      output(30) => mem_array(30)(430),
      output(31) => mem_array(31)(430),
      output(32) => mem_array(32)(430),
      output(33) => mem_array(33)(430),
      output(34) => mem_array(34)(430),
      output(35) => mem_array(35)(430)
      );
  rom431 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(431),
      output(0)  => mem_array(0)(431),
      output(1)  => mem_array(1)(431),
      output(2)  => mem_array(2)(431),
      output(3)  => mem_array(3)(431),
      output(4)  => mem_array(4)(431),
      output(5)  => mem_array(5)(431),
      output(6)  => mem_array(6)(431),
      output(7)  => mem_array(7)(431),
      output(8)  => mem_array(8)(431),
      output(9)  => mem_array(9)(431),
      output(10) => mem_array(10)(431),
      output(11) => mem_array(11)(431),
      output(12) => mem_array(12)(431),
      output(13) => mem_array(13)(431),
      output(14) => mem_array(14)(431),
      output(15) => mem_array(15)(431),
      output(16) => mem_array(16)(431),
      output(17) => mem_array(17)(431),
      output(18) => mem_array(18)(431),
      output(19) => mem_array(19)(431),
      output(20) => mem_array(20)(431),
      output(21) => mem_array(21)(431),
      output(22) => mem_array(22)(431),
      output(23) => mem_array(23)(431),
      output(24) => mem_array(24)(431),
      output(25) => mem_array(25)(431),
      output(26) => mem_array(26)(431),
      output(27) => mem_array(27)(431),
      output(28) => mem_array(28)(431),
      output(29) => mem_array(29)(431),
      output(30) => mem_array(30)(431),
      output(31) => mem_array(31)(431),
      output(32) => mem_array(32)(431),
      output(33) => mem_array(33)(431),
      output(34) => mem_array(34)(431),
      output(35) => mem_array(35)(431)
      );
  rom432 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(432),
      output(0)  => mem_array(0)(432),
      output(1)  => mem_array(1)(432),
      output(2)  => mem_array(2)(432),
      output(3)  => mem_array(3)(432),
      output(4)  => mem_array(4)(432),
      output(5)  => mem_array(5)(432),
      output(6)  => mem_array(6)(432),
      output(7)  => mem_array(7)(432),
      output(8)  => mem_array(8)(432),
      output(9)  => mem_array(9)(432),
      output(10) => mem_array(10)(432),
      output(11) => mem_array(11)(432),
      output(12) => mem_array(12)(432),
      output(13) => mem_array(13)(432),
      output(14) => mem_array(14)(432),
      output(15) => mem_array(15)(432),
      output(16) => mem_array(16)(432),
      output(17) => mem_array(17)(432),
      output(18) => mem_array(18)(432),
      output(19) => mem_array(19)(432),
      output(20) => mem_array(20)(432),
      output(21) => mem_array(21)(432),
      output(22) => mem_array(22)(432),
      output(23) => mem_array(23)(432),
      output(24) => mem_array(24)(432),
      output(25) => mem_array(25)(432),
      output(26) => mem_array(26)(432),
      output(27) => mem_array(27)(432),
      output(28) => mem_array(28)(432),
      output(29) => mem_array(29)(432),
      output(30) => mem_array(30)(432),
      output(31) => mem_array(31)(432),
      output(32) => mem_array(32)(432),
      output(33) => mem_array(33)(432),
      output(34) => mem_array(34)(432),
      output(35) => mem_array(35)(432)
      );
  rom433 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(433),
      output(0)  => mem_array(0)(433),
      output(1)  => mem_array(1)(433),
      output(2)  => mem_array(2)(433),
      output(3)  => mem_array(3)(433),
      output(4)  => mem_array(4)(433),
      output(5)  => mem_array(5)(433),
      output(6)  => mem_array(6)(433),
      output(7)  => mem_array(7)(433),
      output(8)  => mem_array(8)(433),
      output(9)  => mem_array(9)(433),
      output(10) => mem_array(10)(433),
      output(11) => mem_array(11)(433),
      output(12) => mem_array(12)(433),
      output(13) => mem_array(13)(433),
      output(14) => mem_array(14)(433),
      output(15) => mem_array(15)(433),
      output(16) => mem_array(16)(433),
      output(17) => mem_array(17)(433),
      output(18) => mem_array(18)(433),
      output(19) => mem_array(19)(433),
      output(20) => mem_array(20)(433),
      output(21) => mem_array(21)(433),
      output(22) => mem_array(22)(433),
      output(23) => mem_array(23)(433),
      output(24) => mem_array(24)(433),
      output(25) => mem_array(25)(433),
      output(26) => mem_array(26)(433),
      output(27) => mem_array(27)(433),
      output(28) => mem_array(28)(433),
      output(29) => mem_array(29)(433),
      output(30) => mem_array(30)(433),
      output(31) => mem_array(31)(433),
      output(32) => mem_array(32)(433),
      output(33) => mem_array(33)(433),
      output(34) => mem_array(34)(433),
      output(35) => mem_array(35)(433)
      );
  rom434 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(434),
      output(0)  => mem_array(0)(434),
      output(1)  => mem_array(1)(434),
      output(2)  => mem_array(2)(434),
      output(3)  => mem_array(3)(434),
      output(4)  => mem_array(4)(434),
      output(5)  => mem_array(5)(434),
      output(6)  => mem_array(6)(434),
      output(7)  => mem_array(7)(434),
      output(8)  => mem_array(8)(434),
      output(9)  => mem_array(9)(434),
      output(10) => mem_array(10)(434),
      output(11) => mem_array(11)(434),
      output(12) => mem_array(12)(434),
      output(13) => mem_array(13)(434),
      output(14) => mem_array(14)(434),
      output(15) => mem_array(15)(434),
      output(16) => mem_array(16)(434),
      output(17) => mem_array(17)(434),
      output(18) => mem_array(18)(434),
      output(19) => mem_array(19)(434),
      output(20) => mem_array(20)(434),
      output(21) => mem_array(21)(434),
      output(22) => mem_array(22)(434),
      output(23) => mem_array(23)(434),
      output(24) => mem_array(24)(434),
      output(25) => mem_array(25)(434),
      output(26) => mem_array(26)(434),
      output(27) => mem_array(27)(434),
      output(28) => mem_array(28)(434),
      output(29) => mem_array(29)(434),
      output(30) => mem_array(30)(434),
      output(31) => mem_array(31)(434),
      output(32) => mem_array(32)(434),
      output(33) => mem_array(33)(434),
      output(34) => mem_array(34)(434),
      output(35) => mem_array(35)(434)
      );
  rom435 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(435),
      output(0)  => mem_array(0)(435),
      output(1)  => mem_array(1)(435),
      output(2)  => mem_array(2)(435),
      output(3)  => mem_array(3)(435),
      output(4)  => mem_array(4)(435),
      output(5)  => mem_array(5)(435),
      output(6)  => mem_array(6)(435),
      output(7)  => mem_array(7)(435),
      output(8)  => mem_array(8)(435),
      output(9)  => mem_array(9)(435),
      output(10) => mem_array(10)(435),
      output(11) => mem_array(11)(435),
      output(12) => mem_array(12)(435),
      output(13) => mem_array(13)(435),
      output(14) => mem_array(14)(435),
      output(15) => mem_array(15)(435),
      output(16) => mem_array(16)(435),
      output(17) => mem_array(17)(435),
      output(18) => mem_array(18)(435),
      output(19) => mem_array(19)(435),
      output(20) => mem_array(20)(435),
      output(21) => mem_array(21)(435),
      output(22) => mem_array(22)(435),
      output(23) => mem_array(23)(435),
      output(24) => mem_array(24)(435),
      output(25) => mem_array(25)(435),
      output(26) => mem_array(26)(435),
      output(27) => mem_array(27)(435),
      output(28) => mem_array(28)(435),
      output(29) => mem_array(29)(435),
      output(30) => mem_array(30)(435),
      output(31) => mem_array(31)(435),
      output(32) => mem_array(32)(435),
      output(33) => mem_array(33)(435),
      output(34) => mem_array(34)(435),
      output(35) => mem_array(35)(435)
      );
  rom436 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(436),
      output(0)  => mem_array(0)(436),
      output(1)  => mem_array(1)(436),
      output(2)  => mem_array(2)(436),
      output(3)  => mem_array(3)(436),
      output(4)  => mem_array(4)(436),
      output(5)  => mem_array(5)(436),
      output(6)  => mem_array(6)(436),
      output(7)  => mem_array(7)(436),
      output(8)  => mem_array(8)(436),
      output(9)  => mem_array(9)(436),
      output(10) => mem_array(10)(436),
      output(11) => mem_array(11)(436),
      output(12) => mem_array(12)(436),
      output(13) => mem_array(13)(436),
      output(14) => mem_array(14)(436),
      output(15) => mem_array(15)(436),
      output(16) => mem_array(16)(436),
      output(17) => mem_array(17)(436),
      output(18) => mem_array(18)(436),
      output(19) => mem_array(19)(436),
      output(20) => mem_array(20)(436),
      output(21) => mem_array(21)(436),
      output(22) => mem_array(22)(436),
      output(23) => mem_array(23)(436),
      output(24) => mem_array(24)(436),
      output(25) => mem_array(25)(436),
      output(26) => mem_array(26)(436),
      output(27) => mem_array(27)(436),
      output(28) => mem_array(28)(436),
      output(29) => mem_array(29)(436),
      output(30) => mem_array(30)(436),
      output(31) => mem_array(31)(436),
      output(32) => mem_array(32)(436),
      output(33) => mem_array(33)(436),
      output(34) => mem_array(34)(436),
      output(35) => mem_array(35)(436)
      );
  rom437 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(437),
      output(0)  => mem_array(0)(437),
      output(1)  => mem_array(1)(437),
      output(2)  => mem_array(2)(437),
      output(3)  => mem_array(3)(437),
      output(4)  => mem_array(4)(437),
      output(5)  => mem_array(5)(437),
      output(6)  => mem_array(6)(437),
      output(7)  => mem_array(7)(437),
      output(8)  => mem_array(8)(437),
      output(9)  => mem_array(9)(437),
      output(10) => mem_array(10)(437),
      output(11) => mem_array(11)(437),
      output(12) => mem_array(12)(437),
      output(13) => mem_array(13)(437),
      output(14) => mem_array(14)(437),
      output(15) => mem_array(15)(437),
      output(16) => mem_array(16)(437),
      output(17) => mem_array(17)(437),
      output(18) => mem_array(18)(437),
      output(19) => mem_array(19)(437),
      output(20) => mem_array(20)(437),
      output(21) => mem_array(21)(437),
      output(22) => mem_array(22)(437),
      output(23) => mem_array(23)(437),
      output(24) => mem_array(24)(437),
      output(25) => mem_array(25)(437),
      output(26) => mem_array(26)(437),
      output(27) => mem_array(27)(437),
      output(28) => mem_array(28)(437),
      output(29) => mem_array(29)(437),
      output(30) => mem_array(30)(437),
      output(31) => mem_array(31)(437),
      output(32) => mem_array(32)(437),
      output(33) => mem_array(33)(437),
      output(34) => mem_array(34)(437),
      output(35) => mem_array(35)(437)
      );
  rom438 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(438),
      output(0)  => mem_array(0)(438),
      output(1)  => mem_array(1)(438),
      output(2)  => mem_array(2)(438),
      output(3)  => mem_array(3)(438),
      output(4)  => mem_array(4)(438),
      output(5)  => mem_array(5)(438),
      output(6)  => mem_array(6)(438),
      output(7)  => mem_array(7)(438),
      output(8)  => mem_array(8)(438),
      output(9)  => mem_array(9)(438),
      output(10) => mem_array(10)(438),
      output(11) => mem_array(11)(438),
      output(12) => mem_array(12)(438),
      output(13) => mem_array(13)(438),
      output(14) => mem_array(14)(438),
      output(15) => mem_array(15)(438),
      output(16) => mem_array(16)(438),
      output(17) => mem_array(17)(438),
      output(18) => mem_array(18)(438),
      output(19) => mem_array(19)(438),
      output(20) => mem_array(20)(438),
      output(21) => mem_array(21)(438),
      output(22) => mem_array(22)(438),
      output(23) => mem_array(23)(438),
      output(24) => mem_array(24)(438),
      output(25) => mem_array(25)(438),
      output(26) => mem_array(26)(438),
      output(27) => mem_array(27)(438),
      output(28) => mem_array(28)(438),
      output(29) => mem_array(29)(438),
      output(30) => mem_array(30)(438),
      output(31) => mem_array(31)(438),
      output(32) => mem_array(32)(438),
      output(33) => mem_array(33)(438),
      output(34) => mem_array(34)(438),
      output(35) => mem_array(35)(438)
      );
  rom439 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(439),
      output(0)  => mem_array(0)(439),
      output(1)  => mem_array(1)(439),
      output(2)  => mem_array(2)(439),
      output(3)  => mem_array(3)(439),
      output(4)  => mem_array(4)(439),
      output(5)  => mem_array(5)(439),
      output(6)  => mem_array(6)(439),
      output(7)  => mem_array(7)(439),
      output(8)  => mem_array(8)(439),
      output(9)  => mem_array(9)(439),
      output(10) => mem_array(10)(439),
      output(11) => mem_array(11)(439),
      output(12) => mem_array(12)(439),
      output(13) => mem_array(13)(439),
      output(14) => mem_array(14)(439),
      output(15) => mem_array(15)(439),
      output(16) => mem_array(16)(439),
      output(17) => mem_array(17)(439),
      output(18) => mem_array(18)(439),
      output(19) => mem_array(19)(439),
      output(20) => mem_array(20)(439),
      output(21) => mem_array(21)(439),
      output(22) => mem_array(22)(439),
      output(23) => mem_array(23)(439),
      output(24) => mem_array(24)(439),
      output(25) => mem_array(25)(439),
      output(26) => mem_array(26)(439),
      output(27) => mem_array(27)(439),
      output(28) => mem_array(28)(439),
      output(29) => mem_array(29)(439),
      output(30) => mem_array(30)(439),
      output(31) => mem_array(31)(439),
      output(32) => mem_array(32)(439),
      output(33) => mem_array(33)(439),
      output(34) => mem_array(34)(439),
      output(35) => mem_array(35)(439)
      );
  rom440 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(440),
      output(0)  => mem_array(0)(440),
      output(1)  => mem_array(1)(440),
      output(2)  => mem_array(2)(440),
      output(3)  => mem_array(3)(440),
      output(4)  => mem_array(4)(440),
      output(5)  => mem_array(5)(440),
      output(6)  => mem_array(6)(440),
      output(7)  => mem_array(7)(440),
      output(8)  => mem_array(8)(440),
      output(9)  => mem_array(9)(440),
      output(10) => mem_array(10)(440),
      output(11) => mem_array(11)(440),
      output(12) => mem_array(12)(440),
      output(13) => mem_array(13)(440),
      output(14) => mem_array(14)(440),
      output(15) => mem_array(15)(440),
      output(16) => mem_array(16)(440),
      output(17) => mem_array(17)(440),
      output(18) => mem_array(18)(440),
      output(19) => mem_array(19)(440),
      output(20) => mem_array(20)(440),
      output(21) => mem_array(21)(440),
      output(22) => mem_array(22)(440),
      output(23) => mem_array(23)(440),
      output(24) => mem_array(24)(440),
      output(25) => mem_array(25)(440),
      output(26) => mem_array(26)(440),
      output(27) => mem_array(27)(440),
      output(28) => mem_array(28)(440),
      output(29) => mem_array(29)(440),
      output(30) => mem_array(30)(440),
      output(31) => mem_array(31)(440),
      output(32) => mem_array(32)(440),
      output(33) => mem_array(33)(440),
      output(34) => mem_array(34)(440),
      output(35) => mem_array(35)(440)
      );
  rom441 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(441),
      output(0)  => mem_array(0)(441),
      output(1)  => mem_array(1)(441),
      output(2)  => mem_array(2)(441),
      output(3)  => mem_array(3)(441),
      output(4)  => mem_array(4)(441),
      output(5)  => mem_array(5)(441),
      output(6)  => mem_array(6)(441),
      output(7)  => mem_array(7)(441),
      output(8)  => mem_array(8)(441),
      output(9)  => mem_array(9)(441),
      output(10) => mem_array(10)(441),
      output(11) => mem_array(11)(441),
      output(12) => mem_array(12)(441),
      output(13) => mem_array(13)(441),
      output(14) => mem_array(14)(441),
      output(15) => mem_array(15)(441),
      output(16) => mem_array(16)(441),
      output(17) => mem_array(17)(441),
      output(18) => mem_array(18)(441),
      output(19) => mem_array(19)(441),
      output(20) => mem_array(20)(441),
      output(21) => mem_array(21)(441),
      output(22) => mem_array(22)(441),
      output(23) => mem_array(23)(441),
      output(24) => mem_array(24)(441),
      output(25) => mem_array(25)(441),
      output(26) => mem_array(26)(441),
      output(27) => mem_array(27)(441),
      output(28) => mem_array(28)(441),
      output(29) => mem_array(29)(441),
      output(30) => mem_array(30)(441),
      output(31) => mem_array(31)(441),
      output(32) => mem_array(32)(441),
      output(33) => mem_array(33)(441),
      output(34) => mem_array(34)(441),
      output(35) => mem_array(35)(441)
      );
  rom442 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(442),
      output(0)  => mem_array(0)(442),
      output(1)  => mem_array(1)(442),
      output(2)  => mem_array(2)(442),
      output(3)  => mem_array(3)(442),
      output(4)  => mem_array(4)(442),
      output(5)  => mem_array(5)(442),
      output(6)  => mem_array(6)(442),
      output(7)  => mem_array(7)(442),
      output(8)  => mem_array(8)(442),
      output(9)  => mem_array(9)(442),
      output(10) => mem_array(10)(442),
      output(11) => mem_array(11)(442),
      output(12) => mem_array(12)(442),
      output(13) => mem_array(13)(442),
      output(14) => mem_array(14)(442),
      output(15) => mem_array(15)(442),
      output(16) => mem_array(16)(442),
      output(17) => mem_array(17)(442),
      output(18) => mem_array(18)(442),
      output(19) => mem_array(19)(442),
      output(20) => mem_array(20)(442),
      output(21) => mem_array(21)(442),
      output(22) => mem_array(22)(442),
      output(23) => mem_array(23)(442),
      output(24) => mem_array(24)(442),
      output(25) => mem_array(25)(442),
      output(26) => mem_array(26)(442),
      output(27) => mem_array(27)(442),
      output(28) => mem_array(28)(442),
      output(29) => mem_array(29)(442),
      output(30) => mem_array(30)(442),
      output(31) => mem_array(31)(442),
      output(32) => mem_array(32)(442),
      output(33) => mem_array(33)(442),
      output(34) => mem_array(34)(442),
      output(35) => mem_array(35)(442)
      );
  rom443 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(443),
      output(0)  => mem_array(0)(443),
      output(1)  => mem_array(1)(443),
      output(2)  => mem_array(2)(443),
      output(3)  => mem_array(3)(443),
      output(4)  => mem_array(4)(443),
      output(5)  => mem_array(5)(443),
      output(6)  => mem_array(6)(443),
      output(7)  => mem_array(7)(443),
      output(8)  => mem_array(8)(443),
      output(9)  => mem_array(9)(443),
      output(10) => mem_array(10)(443),
      output(11) => mem_array(11)(443),
      output(12) => mem_array(12)(443),
      output(13) => mem_array(13)(443),
      output(14) => mem_array(14)(443),
      output(15) => mem_array(15)(443),
      output(16) => mem_array(16)(443),
      output(17) => mem_array(17)(443),
      output(18) => mem_array(18)(443),
      output(19) => mem_array(19)(443),
      output(20) => mem_array(20)(443),
      output(21) => mem_array(21)(443),
      output(22) => mem_array(22)(443),
      output(23) => mem_array(23)(443),
      output(24) => mem_array(24)(443),
      output(25) => mem_array(25)(443),
      output(26) => mem_array(26)(443),
      output(27) => mem_array(27)(443),
      output(28) => mem_array(28)(443),
      output(29) => mem_array(29)(443),
      output(30) => mem_array(30)(443),
      output(31) => mem_array(31)(443),
      output(32) => mem_array(32)(443),
      output(33) => mem_array(33)(443),
      output(34) => mem_array(34)(443),
      output(35) => mem_array(35)(443)
      );
  rom444 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(444),
      output(0)  => mem_array(0)(444),
      output(1)  => mem_array(1)(444),
      output(2)  => mem_array(2)(444),
      output(3)  => mem_array(3)(444),
      output(4)  => mem_array(4)(444),
      output(5)  => mem_array(5)(444),
      output(6)  => mem_array(6)(444),
      output(7)  => mem_array(7)(444),
      output(8)  => mem_array(8)(444),
      output(9)  => mem_array(9)(444),
      output(10) => mem_array(10)(444),
      output(11) => mem_array(11)(444),
      output(12) => mem_array(12)(444),
      output(13) => mem_array(13)(444),
      output(14) => mem_array(14)(444),
      output(15) => mem_array(15)(444),
      output(16) => mem_array(16)(444),
      output(17) => mem_array(17)(444),
      output(18) => mem_array(18)(444),
      output(19) => mem_array(19)(444),
      output(20) => mem_array(20)(444),
      output(21) => mem_array(21)(444),
      output(22) => mem_array(22)(444),
      output(23) => mem_array(23)(444),
      output(24) => mem_array(24)(444),
      output(25) => mem_array(25)(444),
      output(26) => mem_array(26)(444),
      output(27) => mem_array(27)(444),
      output(28) => mem_array(28)(444),
      output(29) => mem_array(29)(444),
      output(30) => mem_array(30)(444),
      output(31) => mem_array(31)(444),
      output(32) => mem_array(32)(444),
      output(33) => mem_array(33)(444),
      output(34) => mem_array(34)(444),
      output(35) => mem_array(35)(444)
      );
  rom445 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(445),
      output(0)  => mem_array(0)(445),
      output(1)  => mem_array(1)(445),
      output(2)  => mem_array(2)(445),
      output(3)  => mem_array(3)(445),
      output(4)  => mem_array(4)(445),
      output(5)  => mem_array(5)(445),
      output(6)  => mem_array(6)(445),
      output(7)  => mem_array(7)(445),
      output(8)  => mem_array(8)(445),
      output(9)  => mem_array(9)(445),
      output(10) => mem_array(10)(445),
      output(11) => mem_array(11)(445),
      output(12) => mem_array(12)(445),
      output(13) => mem_array(13)(445),
      output(14) => mem_array(14)(445),
      output(15) => mem_array(15)(445),
      output(16) => mem_array(16)(445),
      output(17) => mem_array(17)(445),
      output(18) => mem_array(18)(445),
      output(19) => mem_array(19)(445),
      output(20) => mem_array(20)(445),
      output(21) => mem_array(21)(445),
      output(22) => mem_array(22)(445),
      output(23) => mem_array(23)(445),
      output(24) => mem_array(24)(445),
      output(25) => mem_array(25)(445),
      output(26) => mem_array(26)(445),
      output(27) => mem_array(27)(445),
      output(28) => mem_array(28)(445),
      output(29) => mem_array(29)(445),
      output(30) => mem_array(30)(445),
      output(31) => mem_array(31)(445),
      output(32) => mem_array(32)(445),
      output(33) => mem_array(33)(445),
      output(34) => mem_array(34)(445),
      output(35) => mem_array(35)(445)
      );
  rom446 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(446),
      output(0)  => mem_array(0)(446),
      output(1)  => mem_array(1)(446),
      output(2)  => mem_array(2)(446),
      output(3)  => mem_array(3)(446),
      output(4)  => mem_array(4)(446),
      output(5)  => mem_array(5)(446),
      output(6)  => mem_array(6)(446),
      output(7)  => mem_array(7)(446),
      output(8)  => mem_array(8)(446),
      output(9)  => mem_array(9)(446),
      output(10) => mem_array(10)(446),
      output(11) => mem_array(11)(446),
      output(12) => mem_array(12)(446),
      output(13) => mem_array(13)(446),
      output(14) => mem_array(14)(446),
      output(15) => mem_array(15)(446),
      output(16) => mem_array(16)(446),
      output(17) => mem_array(17)(446),
      output(18) => mem_array(18)(446),
      output(19) => mem_array(19)(446),
      output(20) => mem_array(20)(446),
      output(21) => mem_array(21)(446),
      output(22) => mem_array(22)(446),
      output(23) => mem_array(23)(446),
      output(24) => mem_array(24)(446),
      output(25) => mem_array(25)(446),
      output(26) => mem_array(26)(446),
      output(27) => mem_array(27)(446),
      output(28) => mem_array(28)(446),
      output(29) => mem_array(29)(446),
      output(30) => mem_array(30)(446),
      output(31) => mem_array(31)(446),
      output(32) => mem_array(32)(446),
      output(33) => mem_array(33)(446),
      output(34) => mem_array(34)(446),
      output(35) => mem_array(35)(446)
      );
  rom447 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(447),
      output(0)  => mem_array(0)(447),
      output(1)  => mem_array(1)(447),
      output(2)  => mem_array(2)(447),
      output(3)  => mem_array(3)(447),
      output(4)  => mem_array(4)(447),
      output(5)  => mem_array(5)(447),
      output(6)  => mem_array(6)(447),
      output(7)  => mem_array(7)(447),
      output(8)  => mem_array(8)(447),
      output(9)  => mem_array(9)(447),
      output(10) => mem_array(10)(447),
      output(11) => mem_array(11)(447),
      output(12) => mem_array(12)(447),
      output(13) => mem_array(13)(447),
      output(14) => mem_array(14)(447),
      output(15) => mem_array(15)(447),
      output(16) => mem_array(16)(447),
      output(17) => mem_array(17)(447),
      output(18) => mem_array(18)(447),
      output(19) => mem_array(19)(447),
      output(20) => mem_array(20)(447),
      output(21) => mem_array(21)(447),
      output(22) => mem_array(22)(447),
      output(23) => mem_array(23)(447),
      output(24) => mem_array(24)(447),
      output(25) => mem_array(25)(447),
      output(26) => mem_array(26)(447),
      output(27) => mem_array(27)(447),
      output(28) => mem_array(28)(447),
      output(29) => mem_array(29)(447),
      output(30) => mem_array(30)(447),
      output(31) => mem_array(31)(447),
      output(32) => mem_array(32)(447),
      output(33) => mem_array(33)(447),
      output(34) => mem_array(34)(447),
      output(35) => mem_array(35)(447)
      );
  rom448 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(448),
      output(0)  => mem_array(0)(448),
      output(1)  => mem_array(1)(448),
      output(2)  => mem_array(2)(448),
      output(3)  => mem_array(3)(448),
      output(4)  => mem_array(4)(448),
      output(5)  => mem_array(5)(448),
      output(6)  => mem_array(6)(448),
      output(7)  => mem_array(7)(448),
      output(8)  => mem_array(8)(448),
      output(9)  => mem_array(9)(448),
      output(10) => mem_array(10)(448),
      output(11) => mem_array(11)(448),
      output(12) => mem_array(12)(448),
      output(13) => mem_array(13)(448),
      output(14) => mem_array(14)(448),
      output(15) => mem_array(15)(448),
      output(16) => mem_array(16)(448),
      output(17) => mem_array(17)(448),
      output(18) => mem_array(18)(448),
      output(19) => mem_array(19)(448),
      output(20) => mem_array(20)(448),
      output(21) => mem_array(21)(448),
      output(22) => mem_array(22)(448),
      output(23) => mem_array(23)(448),
      output(24) => mem_array(24)(448),
      output(25) => mem_array(25)(448),
      output(26) => mem_array(26)(448),
      output(27) => mem_array(27)(448),
      output(28) => mem_array(28)(448),
      output(29) => mem_array(29)(448),
      output(30) => mem_array(30)(448),
      output(31) => mem_array(31)(448),
      output(32) => mem_array(32)(448),
      output(33) => mem_array(33)(448),
      output(34) => mem_array(34)(448),
      output(35) => mem_array(35)(448)
      );
  rom449 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(449),
      output(0)  => mem_array(0)(449),
      output(1)  => mem_array(1)(449),
      output(2)  => mem_array(2)(449),
      output(3)  => mem_array(3)(449),
      output(4)  => mem_array(4)(449),
      output(5)  => mem_array(5)(449),
      output(6)  => mem_array(6)(449),
      output(7)  => mem_array(7)(449),
      output(8)  => mem_array(8)(449),
      output(9)  => mem_array(9)(449),
      output(10) => mem_array(10)(449),
      output(11) => mem_array(11)(449),
      output(12) => mem_array(12)(449),
      output(13) => mem_array(13)(449),
      output(14) => mem_array(14)(449),
      output(15) => mem_array(15)(449),
      output(16) => mem_array(16)(449),
      output(17) => mem_array(17)(449),
      output(18) => mem_array(18)(449),
      output(19) => mem_array(19)(449),
      output(20) => mem_array(20)(449),
      output(21) => mem_array(21)(449),
      output(22) => mem_array(22)(449),
      output(23) => mem_array(23)(449),
      output(24) => mem_array(24)(449),
      output(25) => mem_array(25)(449),
      output(26) => mem_array(26)(449),
      output(27) => mem_array(27)(449),
      output(28) => mem_array(28)(449),
      output(29) => mem_array(29)(449),
      output(30) => mem_array(30)(449),
      output(31) => mem_array(31)(449),
      output(32) => mem_array(32)(449),
      output(33) => mem_array(33)(449),
      output(34) => mem_array(34)(449),
      output(35) => mem_array(35)(449)
      );
  rom450 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(450),
      output(0)  => mem_array(0)(450),
      output(1)  => mem_array(1)(450),
      output(2)  => mem_array(2)(450),
      output(3)  => mem_array(3)(450),
      output(4)  => mem_array(4)(450),
      output(5)  => mem_array(5)(450),
      output(6)  => mem_array(6)(450),
      output(7)  => mem_array(7)(450),
      output(8)  => mem_array(8)(450),
      output(9)  => mem_array(9)(450),
      output(10) => mem_array(10)(450),
      output(11) => mem_array(11)(450),
      output(12) => mem_array(12)(450),
      output(13) => mem_array(13)(450),
      output(14) => mem_array(14)(450),
      output(15) => mem_array(15)(450),
      output(16) => mem_array(16)(450),
      output(17) => mem_array(17)(450),
      output(18) => mem_array(18)(450),
      output(19) => mem_array(19)(450),
      output(20) => mem_array(20)(450),
      output(21) => mem_array(21)(450),
      output(22) => mem_array(22)(450),
      output(23) => mem_array(23)(450),
      output(24) => mem_array(24)(450),
      output(25) => mem_array(25)(450),
      output(26) => mem_array(26)(450),
      output(27) => mem_array(27)(450),
      output(28) => mem_array(28)(450),
      output(29) => mem_array(29)(450),
      output(30) => mem_array(30)(450),
      output(31) => mem_array(31)(450),
      output(32) => mem_array(32)(450),
      output(33) => mem_array(33)(450),
      output(34) => mem_array(34)(450),
      output(35) => mem_array(35)(450)
      );
  rom451 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(451),
      output(0)  => mem_array(0)(451),
      output(1)  => mem_array(1)(451),
      output(2)  => mem_array(2)(451),
      output(3)  => mem_array(3)(451),
      output(4)  => mem_array(4)(451),
      output(5)  => mem_array(5)(451),
      output(6)  => mem_array(6)(451),
      output(7)  => mem_array(7)(451),
      output(8)  => mem_array(8)(451),
      output(9)  => mem_array(9)(451),
      output(10) => mem_array(10)(451),
      output(11) => mem_array(11)(451),
      output(12) => mem_array(12)(451),
      output(13) => mem_array(13)(451),
      output(14) => mem_array(14)(451),
      output(15) => mem_array(15)(451),
      output(16) => mem_array(16)(451),
      output(17) => mem_array(17)(451),
      output(18) => mem_array(18)(451),
      output(19) => mem_array(19)(451),
      output(20) => mem_array(20)(451),
      output(21) => mem_array(21)(451),
      output(22) => mem_array(22)(451),
      output(23) => mem_array(23)(451),
      output(24) => mem_array(24)(451),
      output(25) => mem_array(25)(451),
      output(26) => mem_array(26)(451),
      output(27) => mem_array(27)(451),
      output(28) => mem_array(28)(451),
      output(29) => mem_array(29)(451),
      output(30) => mem_array(30)(451),
      output(31) => mem_array(31)(451),
      output(32) => mem_array(32)(451),
      output(33) => mem_array(33)(451),
      output(34) => mem_array(34)(451),
      output(35) => mem_array(35)(451)
      );
  rom452 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(452),
      output(0)  => mem_array(0)(452),
      output(1)  => mem_array(1)(452),
      output(2)  => mem_array(2)(452),
      output(3)  => mem_array(3)(452),
      output(4)  => mem_array(4)(452),
      output(5)  => mem_array(5)(452),
      output(6)  => mem_array(6)(452),
      output(7)  => mem_array(7)(452),
      output(8)  => mem_array(8)(452),
      output(9)  => mem_array(9)(452),
      output(10) => mem_array(10)(452),
      output(11) => mem_array(11)(452),
      output(12) => mem_array(12)(452),
      output(13) => mem_array(13)(452),
      output(14) => mem_array(14)(452),
      output(15) => mem_array(15)(452),
      output(16) => mem_array(16)(452),
      output(17) => mem_array(17)(452),
      output(18) => mem_array(18)(452),
      output(19) => mem_array(19)(452),
      output(20) => mem_array(20)(452),
      output(21) => mem_array(21)(452),
      output(22) => mem_array(22)(452),
      output(23) => mem_array(23)(452),
      output(24) => mem_array(24)(452),
      output(25) => mem_array(25)(452),
      output(26) => mem_array(26)(452),
      output(27) => mem_array(27)(452),
      output(28) => mem_array(28)(452),
      output(29) => mem_array(29)(452),
      output(30) => mem_array(30)(452),
      output(31) => mem_array(31)(452),
      output(32) => mem_array(32)(452),
      output(33) => mem_array(33)(452),
      output(34) => mem_array(34)(452),
      output(35) => mem_array(35)(452)
      );
  rom453 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(453),
      output(0)  => mem_array(0)(453),
      output(1)  => mem_array(1)(453),
      output(2)  => mem_array(2)(453),
      output(3)  => mem_array(3)(453),
      output(4)  => mem_array(4)(453),
      output(5)  => mem_array(5)(453),
      output(6)  => mem_array(6)(453),
      output(7)  => mem_array(7)(453),
      output(8)  => mem_array(8)(453),
      output(9)  => mem_array(9)(453),
      output(10) => mem_array(10)(453),
      output(11) => mem_array(11)(453),
      output(12) => mem_array(12)(453),
      output(13) => mem_array(13)(453),
      output(14) => mem_array(14)(453),
      output(15) => mem_array(15)(453),
      output(16) => mem_array(16)(453),
      output(17) => mem_array(17)(453),
      output(18) => mem_array(18)(453),
      output(19) => mem_array(19)(453),
      output(20) => mem_array(20)(453),
      output(21) => mem_array(21)(453),
      output(22) => mem_array(22)(453),
      output(23) => mem_array(23)(453),
      output(24) => mem_array(24)(453),
      output(25) => mem_array(25)(453),
      output(26) => mem_array(26)(453),
      output(27) => mem_array(27)(453),
      output(28) => mem_array(28)(453),
      output(29) => mem_array(29)(453),
      output(30) => mem_array(30)(453),
      output(31) => mem_array(31)(453),
      output(32) => mem_array(32)(453),
      output(33) => mem_array(33)(453),
      output(34) => mem_array(34)(453),
      output(35) => mem_array(35)(453)
      );
  rom454 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(454),
      output(0)  => mem_array(0)(454),
      output(1)  => mem_array(1)(454),
      output(2)  => mem_array(2)(454),
      output(3)  => mem_array(3)(454),
      output(4)  => mem_array(4)(454),
      output(5)  => mem_array(5)(454),
      output(6)  => mem_array(6)(454),
      output(7)  => mem_array(7)(454),
      output(8)  => mem_array(8)(454),
      output(9)  => mem_array(9)(454),
      output(10) => mem_array(10)(454),
      output(11) => mem_array(11)(454),
      output(12) => mem_array(12)(454),
      output(13) => mem_array(13)(454),
      output(14) => mem_array(14)(454),
      output(15) => mem_array(15)(454),
      output(16) => mem_array(16)(454),
      output(17) => mem_array(17)(454),
      output(18) => mem_array(18)(454),
      output(19) => mem_array(19)(454),
      output(20) => mem_array(20)(454),
      output(21) => mem_array(21)(454),
      output(22) => mem_array(22)(454),
      output(23) => mem_array(23)(454),
      output(24) => mem_array(24)(454),
      output(25) => mem_array(25)(454),
      output(26) => mem_array(26)(454),
      output(27) => mem_array(27)(454),
      output(28) => mem_array(28)(454),
      output(29) => mem_array(29)(454),
      output(30) => mem_array(30)(454),
      output(31) => mem_array(31)(454),
      output(32) => mem_array(32)(454),
      output(33) => mem_array(33)(454),
      output(34) => mem_array(34)(454),
      output(35) => mem_array(35)(454)
      );
  rom455 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(455),
      output(0)  => mem_array(0)(455),
      output(1)  => mem_array(1)(455),
      output(2)  => mem_array(2)(455),
      output(3)  => mem_array(3)(455),
      output(4)  => mem_array(4)(455),
      output(5)  => mem_array(5)(455),
      output(6)  => mem_array(6)(455),
      output(7)  => mem_array(7)(455),
      output(8)  => mem_array(8)(455),
      output(9)  => mem_array(9)(455),
      output(10) => mem_array(10)(455),
      output(11) => mem_array(11)(455),
      output(12) => mem_array(12)(455),
      output(13) => mem_array(13)(455),
      output(14) => mem_array(14)(455),
      output(15) => mem_array(15)(455),
      output(16) => mem_array(16)(455),
      output(17) => mem_array(17)(455),
      output(18) => mem_array(18)(455),
      output(19) => mem_array(19)(455),
      output(20) => mem_array(20)(455),
      output(21) => mem_array(21)(455),
      output(22) => mem_array(22)(455),
      output(23) => mem_array(23)(455),
      output(24) => mem_array(24)(455),
      output(25) => mem_array(25)(455),
      output(26) => mem_array(26)(455),
      output(27) => mem_array(27)(455),
      output(28) => mem_array(28)(455),
      output(29) => mem_array(29)(455),
      output(30) => mem_array(30)(455),
      output(31) => mem_array(31)(455),
      output(32) => mem_array(32)(455),
      output(33) => mem_array(33)(455),
      output(34) => mem_array(34)(455),
      output(35) => mem_array(35)(455)
      );
  rom456 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(456),
      output(0)  => mem_array(0)(456),
      output(1)  => mem_array(1)(456),
      output(2)  => mem_array(2)(456),
      output(3)  => mem_array(3)(456),
      output(4)  => mem_array(4)(456),
      output(5)  => mem_array(5)(456),
      output(6)  => mem_array(6)(456),
      output(7)  => mem_array(7)(456),
      output(8)  => mem_array(8)(456),
      output(9)  => mem_array(9)(456),
      output(10) => mem_array(10)(456),
      output(11) => mem_array(11)(456),
      output(12) => mem_array(12)(456),
      output(13) => mem_array(13)(456),
      output(14) => mem_array(14)(456),
      output(15) => mem_array(15)(456),
      output(16) => mem_array(16)(456),
      output(17) => mem_array(17)(456),
      output(18) => mem_array(18)(456),
      output(19) => mem_array(19)(456),
      output(20) => mem_array(20)(456),
      output(21) => mem_array(21)(456),
      output(22) => mem_array(22)(456),
      output(23) => mem_array(23)(456),
      output(24) => mem_array(24)(456),
      output(25) => mem_array(25)(456),
      output(26) => mem_array(26)(456),
      output(27) => mem_array(27)(456),
      output(28) => mem_array(28)(456),
      output(29) => mem_array(29)(456),
      output(30) => mem_array(30)(456),
      output(31) => mem_array(31)(456),
      output(32) => mem_array(32)(456),
      output(33) => mem_array(33)(456),
      output(34) => mem_array(34)(456),
      output(35) => mem_array(35)(456)
      );
  rom457 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(457),
      output(0)  => mem_array(0)(457),
      output(1)  => mem_array(1)(457),
      output(2)  => mem_array(2)(457),
      output(3)  => mem_array(3)(457),
      output(4)  => mem_array(4)(457),
      output(5)  => mem_array(5)(457),
      output(6)  => mem_array(6)(457),
      output(7)  => mem_array(7)(457),
      output(8)  => mem_array(8)(457),
      output(9)  => mem_array(9)(457),
      output(10) => mem_array(10)(457),
      output(11) => mem_array(11)(457),
      output(12) => mem_array(12)(457),
      output(13) => mem_array(13)(457),
      output(14) => mem_array(14)(457),
      output(15) => mem_array(15)(457),
      output(16) => mem_array(16)(457),
      output(17) => mem_array(17)(457),
      output(18) => mem_array(18)(457),
      output(19) => mem_array(19)(457),
      output(20) => mem_array(20)(457),
      output(21) => mem_array(21)(457),
      output(22) => mem_array(22)(457),
      output(23) => mem_array(23)(457),
      output(24) => mem_array(24)(457),
      output(25) => mem_array(25)(457),
      output(26) => mem_array(26)(457),
      output(27) => mem_array(27)(457),
      output(28) => mem_array(28)(457),
      output(29) => mem_array(29)(457),
      output(30) => mem_array(30)(457),
      output(31) => mem_array(31)(457),
      output(32) => mem_array(32)(457),
      output(33) => mem_array(33)(457),
      output(34) => mem_array(34)(457),
      output(35) => mem_array(35)(457)
      );
  rom458 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(458),
      output(0)  => mem_array(0)(458),
      output(1)  => mem_array(1)(458),
      output(2)  => mem_array(2)(458),
      output(3)  => mem_array(3)(458),
      output(4)  => mem_array(4)(458),
      output(5)  => mem_array(5)(458),
      output(6)  => mem_array(6)(458),
      output(7)  => mem_array(7)(458),
      output(8)  => mem_array(8)(458),
      output(9)  => mem_array(9)(458),
      output(10) => mem_array(10)(458),
      output(11) => mem_array(11)(458),
      output(12) => mem_array(12)(458),
      output(13) => mem_array(13)(458),
      output(14) => mem_array(14)(458),
      output(15) => mem_array(15)(458),
      output(16) => mem_array(16)(458),
      output(17) => mem_array(17)(458),
      output(18) => mem_array(18)(458),
      output(19) => mem_array(19)(458),
      output(20) => mem_array(20)(458),
      output(21) => mem_array(21)(458),
      output(22) => mem_array(22)(458),
      output(23) => mem_array(23)(458),
      output(24) => mem_array(24)(458),
      output(25) => mem_array(25)(458),
      output(26) => mem_array(26)(458),
      output(27) => mem_array(27)(458),
      output(28) => mem_array(28)(458),
      output(29) => mem_array(29)(458),
      output(30) => mem_array(30)(458),
      output(31) => mem_array(31)(458),
      output(32) => mem_array(32)(458),
      output(33) => mem_array(33)(458),
      output(34) => mem_array(34)(458),
      output(35) => mem_array(35)(458)
      );
  rom459 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(459),
      output(0)  => mem_array(0)(459),
      output(1)  => mem_array(1)(459),
      output(2)  => mem_array(2)(459),
      output(3)  => mem_array(3)(459),
      output(4)  => mem_array(4)(459),
      output(5)  => mem_array(5)(459),
      output(6)  => mem_array(6)(459),
      output(7)  => mem_array(7)(459),
      output(8)  => mem_array(8)(459),
      output(9)  => mem_array(9)(459),
      output(10) => mem_array(10)(459),
      output(11) => mem_array(11)(459),
      output(12) => mem_array(12)(459),
      output(13) => mem_array(13)(459),
      output(14) => mem_array(14)(459),
      output(15) => mem_array(15)(459),
      output(16) => mem_array(16)(459),
      output(17) => mem_array(17)(459),
      output(18) => mem_array(18)(459),
      output(19) => mem_array(19)(459),
      output(20) => mem_array(20)(459),
      output(21) => mem_array(21)(459),
      output(22) => mem_array(22)(459),
      output(23) => mem_array(23)(459),
      output(24) => mem_array(24)(459),
      output(25) => mem_array(25)(459),
      output(26) => mem_array(26)(459),
      output(27) => mem_array(27)(459),
      output(28) => mem_array(28)(459),
      output(29) => mem_array(29)(459),
      output(30) => mem_array(30)(459),
      output(31) => mem_array(31)(459),
      output(32) => mem_array(32)(459),
      output(33) => mem_array(33)(459),
      output(34) => mem_array(34)(459),
      output(35) => mem_array(35)(459)
      );
  rom460 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(460),
      output(0)  => mem_array(0)(460),
      output(1)  => mem_array(1)(460),
      output(2)  => mem_array(2)(460),
      output(3)  => mem_array(3)(460),
      output(4)  => mem_array(4)(460),
      output(5)  => mem_array(5)(460),
      output(6)  => mem_array(6)(460),
      output(7)  => mem_array(7)(460),
      output(8)  => mem_array(8)(460),
      output(9)  => mem_array(9)(460),
      output(10) => mem_array(10)(460),
      output(11) => mem_array(11)(460),
      output(12) => mem_array(12)(460),
      output(13) => mem_array(13)(460),
      output(14) => mem_array(14)(460),
      output(15) => mem_array(15)(460),
      output(16) => mem_array(16)(460),
      output(17) => mem_array(17)(460),
      output(18) => mem_array(18)(460),
      output(19) => mem_array(19)(460),
      output(20) => mem_array(20)(460),
      output(21) => mem_array(21)(460),
      output(22) => mem_array(22)(460),
      output(23) => mem_array(23)(460),
      output(24) => mem_array(24)(460),
      output(25) => mem_array(25)(460),
      output(26) => mem_array(26)(460),
      output(27) => mem_array(27)(460),
      output(28) => mem_array(28)(460),
      output(29) => mem_array(29)(460),
      output(30) => mem_array(30)(460),
      output(31) => mem_array(31)(460),
      output(32) => mem_array(32)(460),
      output(33) => mem_array(33)(460),
      output(34) => mem_array(34)(460),
      output(35) => mem_array(35)(460)
      );
  rom461 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(461),
      output(0)  => mem_array(0)(461),
      output(1)  => mem_array(1)(461),
      output(2)  => mem_array(2)(461),
      output(3)  => mem_array(3)(461),
      output(4)  => mem_array(4)(461),
      output(5)  => mem_array(5)(461),
      output(6)  => mem_array(6)(461),
      output(7)  => mem_array(7)(461),
      output(8)  => mem_array(8)(461),
      output(9)  => mem_array(9)(461),
      output(10) => mem_array(10)(461),
      output(11) => mem_array(11)(461),
      output(12) => mem_array(12)(461),
      output(13) => mem_array(13)(461),
      output(14) => mem_array(14)(461),
      output(15) => mem_array(15)(461),
      output(16) => mem_array(16)(461),
      output(17) => mem_array(17)(461),
      output(18) => mem_array(18)(461),
      output(19) => mem_array(19)(461),
      output(20) => mem_array(20)(461),
      output(21) => mem_array(21)(461),
      output(22) => mem_array(22)(461),
      output(23) => mem_array(23)(461),
      output(24) => mem_array(24)(461),
      output(25) => mem_array(25)(461),
      output(26) => mem_array(26)(461),
      output(27) => mem_array(27)(461),
      output(28) => mem_array(28)(461),
      output(29) => mem_array(29)(461),
      output(30) => mem_array(30)(461),
      output(31) => mem_array(31)(461),
      output(32) => mem_array(32)(461),
      output(33) => mem_array(33)(461),
      output(34) => mem_array(34)(461),
      output(35) => mem_array(35)(461)
      );
  rom462 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(462),
      output(0)  => mem_array(0)(462),
      output(1)  => mem_array(1)(462),
      output(2)  => mem_array(2)(462),
      output(3)  => mem_array(3)(462),
      output(4)  => mem_array(4)(462),
      output(5)  => mem_array(5)(462),
      output(6)  => mem_array(6)(462),
      output(7)  => mem_array(7)(462),
      output(8)  => mem_array(8)(462),
      output(9)  => mem_array(9)(462),
      output(10) => mem_array(10)(462),
      output(11) => mem_array(11)(462),
      output(12) => mem_array(12)(462),
      output(13) => mem_array(13)(462),
      output(14) => mem_array(14)(462),
      output(15) => mem_array(15)(462),
      output(16) => mem_array(16)(462),
      output(17) => mem_array(17)(462),
      output(18) => mem_array(18)(462),
      output(19) => mem_array(19)(462),
      output(20) => mem_array(20)(462),
      output(21) => mem_array(21)(462),
      output(22) => mem_array(22)(462),
      output(23) => mem_array(23)(462),
      output(24) => mem_array(24)(462),
      output(25) => mem_array(25)(462),
      output(26) => mem_array(26)(462),
      output(27) => mem_array(27)(462),
      output(28) => mem_array(28)(462),
      output(29) => mem_array(29)(462),
      output(30) => mem_array(30)(462),
      output(31) => mem_array(31)(462),
      output(32) => mem_array(32)(462),
      output(33) => mem_array(33)(462),
      output(34) => mem_array(34)(462),
      output(35) => mem_array(35)(462)
      );
  rom463 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(463),
      output(0)  => mem_array(0)(463),
      output(1)  => mem_array(1)(463),
      output(2)  => mem_array(2)(463),
      output(3)  => mem_array(3)(463),
      output(4)  => mem_array(4)(463),
      output(5)  => mem_array(5)(463),
      output(6)  => mem_array(6)(463),
      output(7)  => mem_array(7)(463),
      output(8)  => mem_array(8)(463),
      output(9)  => mem_array(9)(463),
      output(10) => mem_array(10)(463),
      output(11) => mem_array(11)(463),
      output(12) => mem_array(12)(463),
      output(13) => mem_array(13)(463),
      output(14) => mem_array(14)(463),
      output(15) => mem_array(15)(463),
      output(16) => mem_array(16)(463),
      output(17) => mem_array(17)(463),
      output(18) => mem_array(18)(463),
      output(19) => mem_array(19)(463),
      output(20) => mem_array(20)(463),
      output(21) => mem_array(21)(463),
      output(22) => mem_array(22)(463),
      output(23) => mem_array(23)(463),
      output(24) => mem_array(24)(463),
      output(25) => mem_array(25)(463),
      output(26) => mem_array(26)(463),
      output(27) => mem_array(27)(463),
      output(28) => mem_array(28)(463),
      output(29) => mem_array(29)(463),
      output(30) => mem_array(30)(463),
      output(31) => mem_array(31)(463),
      output(32) => mem_array(32)(463),
      output(33) => mem_array(33)(463),
      output(34) => mem_array(34)(463),
      output(35) => mem_array(35)(463)
      );
  rom464 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(464),
      output(0)  => mem_array(0)(464),
      output(1)  => mem_array(1)(464),
      output(2)  => mem_array(2)(464),
      output(3)  => mem_array(3)(464),
      output(4)  => mem_array(4)(464),
      output(5)  => mem_array(5)(464),
      output(6)  => mem_array(6)(464),
      output(7)  => mem_array(7)(464),
      output(8)  => mem_array(8)(464),
      output(9)  => mem_array(9)(464),
      output(10) => mem_array(10)(464),
      output(11) => mem_array(11)(464),
      output(12) => mem_array(12)(464),
      output(13) => mem_array(13)(464),
      output(14) => mem_array(14)(464),
      output(15) => mem_array(15)(464),
      output(16) => mem_array(16)(464),
      output(17) => mem_array(17)(464),
      output(18) => mem_array(18)(464),
      output(19) => mem_array(19)(464),
      output(20) => mem_array(20)(464),
      output(21) => mem_array(21)(464),
      output(22) => mem_array(22)(464),
      output(23) => mem_array(23)(464),
      output(24) => mem_array(24)(464),
      output(25) => mem_array(25)(464),
      output(26) => mem_array(26)(464),
      output(27) => mem_array(27)(464),
      output(28) => mem_array(28)(464),
      output(29) => mem_array(29)(464),
      output(30) => mem_array(30)(464),
      output(31) => mem_array(31)(464),
      output(32) => mem_array(32)(464),
      output(33) => mem_array(33)(464),
      output(34) => mem_array(34)(464),
      output(35) => mem_array(35)(464)
      );
  rom465 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(465),
      output(0)  => mem_array(0)(465),
      output(1)  => mem_array(1)(465),
      output(2)  => mem_array(2)(465),
      output(3)  => mem_array(3)(465),
      output(4)  => mem_array(4)(465),
      output(5)  => mem_array(5)(465),
      output(6)  => mem_array(6)(465),
      output(7)  => mem_array(7)(465),
      output(8)  => mem_array(8)(465),
      output(9)  => mem_array(9)(465),
      output(10) => mem_array(10)(465),
      output(11) => mem_array(11)(465),
      output(12) => mem_array(12)(465),
      output(13) => mem_array(13)(465),
      output(14) => mem_array(14)(465),
      output(15) => mem_array(15)(465),
      output(16) => mem_array(16)(465),
      output(17) => mem_array(17)(465),
      output(18) => mem_array(18)(465),
      output(19) => mem_array(19)(465),
      output(20) => mem_array(20)(465),
      output(21) => mem_array(21)(465),
      output(22) => mem_array(22)(465),
      output(23) => mem_array(23)(465),
      output(24) => mem_array(24)(465),
      output(25) => mem_array(25)(465),
      output(26) => mem_array(26)(465),
      output(27) => mem_array(27)(465),
      output(28) => mem_array(28)(465),
      output(29) => mem_array(29)(465),
      output(30) => mem_array(30)(465),
      output(31) => mem_array(31)(465),
      output(32) => mem_array(32)(465),
      output(33) => mem_array(33)(465),
      output(34) => mem_array(34)(465),
      output(35) => mem_array(35)(465)
      );
  rom466 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(466),
      output(0)  => mem_array(0)(466),
      output(1)  => mem_array(1)(466),
      output(2)  => mem_array(2)(466),
      output(3)  => mem_array(3)(466),
      output(4)  => mem_array(4)(466),
      output(5)  => mem_array(5)(466),
      output(6)  => mem_array(6)(466),
      output(7)  => mem_array(7)(466),
      output(8)  => mem_array(8)(466),
      output(9)  => mem_array(9)(466),
      output(10) => mem_array(10)(466),
      output(11) => mem_array(11)(466),
      output(12) => mem_array(12)(466),
      output(13) => mem_array(13)(466),
      output(14) => mem_array(14)(466),
      output(15) => mem_array(15)(466),
      output(16) => mem_array(16)(466),
      output(17) => mem_array(17)(466),
      output(18) => mem_array(18)(466),
      output(19) => mem_array(19)(466),
      output(20) => mem_array(20)(466),
      output(21) => mem_array(21)(466),
      output(22) => mem_array(22)(466),
      output(23) => mem_array(23)(466),
      output(24) => mem_array(24)(466),
      output(25) => mem_array(25)(466),
      output(26) => mem_array(26)(466),
      output(27) => mem_array(27)(466),
      output(28) => mem_array(28)(466),
      output(29) => mem_array(29)(466),
      output(30) => mem_array(30)(466),
      output(31) => mem_array(31)(466),
      output(32) => mem_array(32)(466),
      output(33) => mem_array(33)(466),
      output(34) => mem_array(34)(466),
      output(35) => mem_array(35)(466)
      );
  rom467 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(467),
      output(0)  => mem_array(0)(467),
      output(1)  => mem_array(1)(467),
      output(2)  => mem_array(2)(467),
      output(3)  => mem_array(3)(467),
      output(4)  => mem_array(4)(467),
      output(5)  => mem_array(5)(467),
      output(6)  => mem_array(6)(467),
      output(7)  => mem_array(7)(467),
      output(8)  => mem_array(8)(467),
      output(9)  => mem_array(9)(467),
      output(10) => mem_array(10)(467),
      output(11) => mem_array(11)(467),
      output(12) => mem_array(12)(467),
      output(13) => mem_array(13)(467),
      output(14) => mem_array(14)(467),
      output(15) => mem_array(15)(467),
      output(16) => mem_array(16)(467),
      output(17) => mem_array(17)(467),
      output(18) => mem_array(18)(467),
      output(19) => mem_array(19)(467),
      output(20) => mem_array(20)(467),
      output(21) => mem_array(21)(467),
      output(22) => mem_array(22)(467),
      output(23) => mem_array(23)(467),
      output(24) => mem_array(24)(467),
      output(25) => mem_array(25)(467),
      output(26) => mem_array(26)(467),
      output(27) => mem_array(27)(467),
      output(28) => mem_array(28)(467),
      output(29) => mem_array(29)(467),
      output(30) => mem_array(30)(467),
      output(31) => mem_array(31)(467),
      output(32) => mem_array(32)(467),
      output(33) => mem_array(33)(467),
      output(34) => mem_array(34)(467),
      output(35) => mem_array(35)(467)
      );
  rom468 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(468),
      output(0)  => mem_array(0)(468),
      output(1)  => mem_array(1)(468),
      output(2)  => mem_array(2)(468),
      output(3)  => mem_array(3)(468),
      output(4)  => mem_array(4)(468),
      output(5)  => mem_array(5)(468),
      output(6)  => mem_array(6)(468),
      output(7)  => mem_array(7)(468),
      output(8)  => mem_array(8)(468),
      output(9)  => mem_array(9)(468),
      output(10) => mem_array(10)(468),
      output(11) => mem_array(11)(468),
      output(12) => mem_array(12)(468),
      output(13) => mem_array(13)(468),
      output(14) => mem_array(14)(468),
      output(15) => mem_array(15)(468),
      output(16) => mem_array(16)(468),
      output(17) => mem_array(17)(468),
      output(18) => mem_array(18)(468),
      output(19) => mem_array(19)(468),
      output(20) => mem_array(20)(468),
      output(21) => mem_array(21)(468),
      output(22) => mem_array(22)(468),
      output(23) => mem_array(23)(468),
      output(24) => mem_array(24)(468),
      output(25) => mem_array(25)(468),
      output(26) => mem_array(26)(468),
      output(27) => mem_array(27)(468),
      output(28) => mem_array(28)(468),
      output(29) => mem_array(29)(468),
      output(30) => mem_array(30)(468),
      output(31) => mem_array(31)(468),
      output(32) => mem_array(32)(468),
      output(33) => mem_array(33)(468),
      output(34) => mem_array(34)(468),
      output(35) => mem_array(35)(468)
      );
  rom469 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(469),
      output(0)  => mem_array(0)(469),
      output(1)  => mem_array(1)(469),
      output(2)  => mem_array(2)(469),
      output(3)  => mem_array(3)(469),
      output(4)  => mem_array(4)(469),
      output(5)  => mem_array(5)(469),
      output(6)  => mem_array(6)(469),
      output(7)  => mem_array(7)(469),
      output(8)  => mem_array(8)(469),
      output(9)  => mem_array(9)(469),
      output(10) => mem_array(10)(469),
      output(11) => mem_array(11)(469),
      output(12) => mem_array(12)(469),
      output(13) => mem_array(13)(469),
      output(14) => mem_array(14)(469),
      output(15) => mem_array(15)(469),
      output(16) => mem_array(16)(469),
      output(17) => mem_array(17)(469),
      output(18) => mem_array(18)(469),
      output(19) => mem_array(19)(469),
      output(20) => mem_array(20)(469),
      output(21) => mem_array(21)(469),
      output(22) => mem_array(22)(469),
      output(23) => mem_array(23)(469),
      output(24) => mem_array(24)(469),
      output(25) => mem_array(25)(469),
      output(26) => mem_array(26)(469),
      output(27) => mem_array(27)(469),
      output(28) => mem_array(28)(469),
      output(29) => mem_array(29)(469),
      output(30) => mem_array(30)(469),
      output(31) => mem_array(31)(469),
      output(32) => mem_array(32)(469),
      output(33) => mem_array(33)(469),
      output(34) => mem_array(34)(469),
      output(35) => mem_array(35)(469)
      );
  rom470 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(470),
      output(0)  => mem_array(0)(470),
      output(1)  => mem_array(1)(470),
      output(2)  => mem_array(2)(470),
      output(3)  => mem_array(3)(470),
      output(4)  => mem_array(4)(470),
      output(5)  => mem_array(5)(470),
      output(6)  => mem_array(6)(470),
      output(7)  => mem_array(7)(470),
      output(8)  => mem_array(8)(470),
      output(9)  => mem_array(9)(470),
      output(10) => mem_array(10)(470),
      output(11) => mem_array(11)(470),
      output(12) => mem_array(12)(470),
      output(13) => mem_array(13)(470),
      output(14) => mem_array(14)(470),
      output(15) => mem_array(15)(470),
      output(16) => mem_array(16)(470),
      output(17) => mem_array(17)(470),
      output(18) => mem_array(18)(470),
      output(19) => mem_array(19)(470),
      output(20) => mem_array(20)(470),
      output(21) => mem_array(21)(470),
      output(22) => mem_array(22)(470),
      output(23) => mem_array(23)(470),
      output(24) => mem_array(24)(470),
      output(25) => mem_array(25)(470),
      output(26) => mem_array(26)(470),
      output(27) => mem_array(27)(470),
      output(28) => mem_array(28)(470),
      output(29) => mem_array(29)(470),
      output(30) => mem_array(30)(470),
      output(31) => mem_array(31)(470),
      output(32) => mem_array(32)(470),
      output(33) => mem_array(33)(470),
      output(34) => mem_array(34)(470),
      output(35) => mem_array(35)(470)
      );
  rom471 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(471),
      output(0)  => mem_array(0)(471),
      output(1)  => mem_array(1)(471),
      output(2)  => mem_array(2)(471),
      output(3)  => mem_array(3)(471),
      output(4)  => mem_array(4)(471),
      output(5)  => mem_array(5)(471),
      output(6)  => mem_array(6)(471),
      output(7)  => mem_array(7)(471),
      output(8)  => mem_array(8)(471),
      output(9)  => mem_array(9)(471),
      output(10) => mem_array(10)(471),
      output(11) => mem_array(11)(471),
      output(12) => mem_array(12)(471),
      output(13) => mem_array(13)(471),
      output(14) => mem_array(14)(471),
      output(15) => mem_array(15)(471),
      output(16) => mem_array(16)(471),
      output(17) => mem_array(17)(471),
      output(18) => mem_array(18)(471),
      output(19) => mem_array(19)(471),
      output(20) => mem_array(20)(471),
      output(21) => mem_array(21)(471),
      output(22) => mem_array(22)(471),
      output(23) => mem_array(23)(471),
      output(24) => mem_array(24)(471),
      output(25) => mem_array(25)(471),
      output(26) => mem_array(26)(471),
      output(27) => mem_array(27)(471),
      output(28) => mem_array(28)(471),
      output(29) => mem_array(29)(471),
      output(30) => mem_array(30)(471),
      output(31) => mem_array(31)(471),
      output(32) => mem_array(32)(471),
      output(33) => mem_array(33)(471),
      output(34) => mem_array(34)(471),
      output(35) => mem_array(35)(471)
      );
  rom472 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(472),
      output(0)  => mem_array(0)(472),
      output(1)  => mem_array(1)(472),
      output(2)  => mem_array(2)(472),
      output(3)  => mem_array(3)(472),
      output(4)  => mem_array(4)(472),
      output(5)  => mem_array(5)(472),
      output(6)  => mem_array(6)(472),
      output(7)  => mem_array(7)(472),
      output(8)  => mem_array(8)(472),
      output(9)  => mem_array(9)(472),
      output(10) => mem_array(10)(472),
      output(11) => mem_array(11)(472),
      output(12) => mem_array(12)(472),
      output(13) => mem_array(13)(472),
      output(14) => mem_array(14)(472),
      output(15) => mem_array(15)(472),
      output(16) => mem_array(16)(472),
      output(17) => mem_array(17)(472),
      output(18) => mem_array(18)(472),
      output(19) => mem_array(19)(472),
      output(20) => mem_array(20)(472),
      output(21) => mem_array(21)(472),
      output(22) => mem_array(22)(472),
      output(23) => mem_array(23)(472),
      output(24) => mem_array(24)(472),
      output(25) => mem_array(25)(472),
      output(26) => mem_array(26)(472),
      output(27) => mem_array(27)(472),
      output(28) => mem_array(28)(472),
      output(29) => mem_array(29)(472),
      output(30) => mem_array(30)(472),
      output(31) => mem_array(31)(472),
      output(32) => mem_array(32)(472),
      output(33) => mem_array(33)(472),
      output(34) => mem_array(34)(472),
      output(35) => mem_array(35)(472)
      );
  rom473 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(473),
      output(0)  => mem_array(0)(473),
      output(1)  => mem_array(1)(473),
      output(2)  => mem_array(2)(473),
      output(3)  => mem_array(3)(473),
      output(4)  => mem_array(4)(473),
      output(5)  => mem_array(5)(473),
      output(6)  => mem_array(6)(473),
      output(7)  => mem_array(7)(473),
      output(8)  => mem_array(8)(473),
      output(9)  => mem_array(9)(473),
      output(10) => mem_array(10)(473),
      output(11) => mem_array(11)(473),
      output(12) => mem_array(12)(473),
      output(13) => mem_array(13)(473),
      output(14) => mem_array(14)(473),
      output(15) => mem_array(15)(473),
      output(16) => mem_array(16)(473),
      output(17) => mem_array(17)(473),
      output(18) => mem_array(18)(473),
      output(19) => mem_array(19)(473),
      output(20) => mem_array(20)(473),
      output(21) => mem_array(21)(473),
      output(22) => mem_array(22)(473),
      output(23) => mem_array(23)(473),
      output(24) => mem_array(24)(473),
      output(25) => mem_array(25)(473),
      output(26) => mem_array(26)(473),
      output(27) => mem_array(27)(473),
      output(28) => mem_array(28)(473),
      output(29) => mem_array(29)(473),
      output(30) => mem_array(30)(473),
      output(31) => mem_array(31)(473),
      output(32) => mem_array(32)(473),
      output(33) => mem_array(33)(473),
      output(34) => mem_array(34)(473),
      output(35) => mem_array(35)(473)
      );
  rom474 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(474),
      output(0)  => mem_array(0)(474),
      output(1)  => mem_array(1)(474),
      output(2)  => mem_array(2)(474),
      output(3)  => mem_array(3)(474),
      output(4)  => mem_array(4)(474),
      output(5)  => mem_array(5)(474),
      output(6)  => mem_array(6)(474),
      output(7)  => mem_array(7)(474),
      output(8)  => mem_array(8)(474),
      output(9)  => mem_array(9)(474),
      output(10) => mem_array(10)(474),
      output(11) => mem_array(11)(474),
      output(12) => mem_array(12)(474),
      output(13) => mem_array(13)(474),
      output(14) => mem_array(14)(474),
      output(15) => mem_array(15)(474),
      output(16) => mem_array(16)(474),
      output(17) => mem_array(17)(474),
      output(18) => mem_array(18)(474),
      output(19) => mem_array(19)(474),
      output(20) => mem_array(20)(474),
      output(21) => mem_array(21)(474),
      output(22) => mem_array(22)(474),
      output(23) => mem_array(23)(474),
      output(24) => mem_array(24)(474),
      output(25) => mem_array(25)(474),
      output(26) => mem_array(26)(474),
      output(27) => mem_array(27)(474),
      output(28) => mem_array(28)(474),
      output(29) => mem_array(29)(474),
      output(30) => mem_array(30)(474),
      output(31) => mem_array(31)(474),
      output(32) => mem_array(32)(474),
      output(33) => mem_array(33)(474),
      output(34) => mem_array(34)(474),
      output(35) => mem_array(35)(474)
      );
  rom475 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(475),
      output(0)  => mem_array(0)(475),
      output(1)  => mem_array(1)(475),
      output(2)  => mem_array(2)(475),
      output(3)  => mem_array(3)(475),
      output(4)  => mem_array(4)(475),
      output(5)  => mem_array(5)(475),
      output(6)  => mem_array(6)(475),
      output(7)  => mem_array(7)(475),
      output(8)  => mem_array(8)(475),
      output(9)  => mem_array(9)(475),
      output(10) => mem_array(10)(475),
      output(11) => mem_array(11)(475),
      output(12) => mem_array(12)(475),
      output(13) => mem_array(13)(475),
      output(14) => mem_array(14)(475),
      output(15) => mem_array(15)(475),
      output(16) => mem_array(16)(475),
      output(17) => mem_array(17)(475),
      output(18) => mem_array(18)(475),
      output(19) => mem_array(19)(475),
      output(20) => mem_array(20)(475),
      output(21) => mem_array(21)(475),
      output(22) => mem_array(22)(475),
      output(23) => mem_array(23)(475),
      output(24) => mem_array(24)(475),
      output(25) => mem_array(25)(475),
      output(26) => mem_array(26)(475),
      output(27) => mem_array(27)(475),
      output(28) => mem_array(28)(475),
      output(29) => mem_array(29)(475),
      output(30) => mem_array(30)(475),
      output(31) => mem_array(31)(475),
      output(32) => mem_array(32)(475),
      output(33) => mem_array(33)(475),
      output(34) => mem_array(34)(475),
      output(35) => mem_array(35)(475)
      );
  rom476 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(476),
      output(0)  => mem_array(0)(476),
      output(1)  => mem_array(1)(476),
      output(2)  => mem_array(2)(476),
      output(3)  => mem_array(3)(476),
      output(4)  => mem_array(4)(476),
      output(5)  => mem_array(5)(476),
      output(6)  => mem_array(6)(476),
      output(7)  => mem_array(7)(476),
      output(8)  => mem_array(8)(476),
      output(9)  => mem_array(9)(476),
      output(10) => mem_array(10)(476),
      output(11) => mem_array(11)(476),
      output(12) => mem_array(12)(476),
      output(13) => mem_array(13)(476),
      output(14) => mem_array(14)(476),
      output(15) => mem_array(15)(476),
      output(16) => mem_array(16)(476),
      output(17) => mem_array(17)(476),
      output(18) => mem_array(18)(476),
      output(19) => mem_array(19)(476),
      output(20) => mem_array(20)(476),
      output(21) => mem_array(21)(476),
      output(22) => mem_array(22)(476),
      output(23) => mem_array(23)(476),
      output(24) => mem_array(24)(476),
      output(25) => mem_array(25)(476),
      output(26) => mem_array(26)(476),
      output(27) => mem_array(27)(476),
      output(28) => mem_array(28)(476),
      output(29) => mem_array(29)(476),
      output(30) => mem_array(30)(476),
      output(31) => mem_array(31)(476),
      output(32) => mem_array(32)(476),
      output(33) => mem_array(33)(476),
      output(34) => mem_array(34)(476),
      output(35) => mem_array(35)(476)
      );
  rom477 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(477),
      output(0)  => mem_array(0)(477),
      output(1)  => mem_array(1)(477),
      output(2)  => mem_array(2)(477),
      output(3)  => mem_array(3)(477),
      output(4)  => mem_array(4)(477),
      output(5)  => mem_array(5)(477),
      output(6)  => mem_array(6)(477),
      output(7)  => mem_array(7)(477),
      output(8)  => mem_array(8)(477),
      output(9)  => mem_array(9)(477),
      output(10) => mem_array(10)(477),
      output(11) => mem_array(11)(477),
      output(12) => mem_array(12)(477),
      output(13) => mem_array(13)(477),
      output(14) => mem_array(14)(477),
      output(15) => mem_array(15)(477),
      output(16) => mem_array(16)(477),
      output(17) => mem_array(17)(477),
      output(18) => mem_array(18)(477),
      output(19) => mem_array(19)(477),
      output(20) => mem_array(20)(477),
      output(21) => mem_array(21)(477),
      output(22) => mem_array(22)(477),
      output(23) => mem_array(23)(477),
      output(24) => mem_array(24)(477),
      output(25) => mem_array(25)(477),
      output(26) => mem_array(26)(477),
      output(27) => mem_array(27)(477),
      output(28) => mem_array(28)(477),
      output(29) => mem_array(29)(477),
      output(30) => mem_array(30)(477),
      output(31) => mem_array(31)(477),
      output(32) => mem_array(32)(477),
      output(33) => mem_array(33)(477),
      output(34) => mem_array(34)(477),
      output(35) => mem_array(35)(477)
      );
  rom478 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(478),
      output(0)  => mem_array(0)(478),
      output(1)  => mem_array(1)(478),
      output(2)  => mem_array(2)(478),
      output(3)  => mem_array(3)(478),
      output(4)  => mem_array(4)(478),
      output(5)  => mem_array(5)(478),
      output(6)  => mem_array(6)(478),
      output(7)  => mem_array(7)(478),
      output(8)  => mem_array(8)(478),
      output(9)  => mem_array(9)(478),
      output(10) => mem_array(10)(478),
      output(11) => mem_array(11)(478),
      output(12) => mem_array(12)(478),
      output(13) => mem_array(13)(478),
      output(14) => mem_array(14)(478),
      output(15) => mem_array(15)(478),
      output(16) => mem_array(16)(478),
      output(17) => mem_array(17)(478),
      output(18) => mem_array(18)(478),
      output(19) => mem_array(19)(478),
      output(20) => mem_array(20)(478),
      output(21) => mem_array(21)(478),
      output(22) => mem_array(22)(478),
      output(23) => mem_array(23)(478),
      output(24) => mem_array(24)(478),
      output(25) => mem_array(25)(478),
      output(26) => mem_array(26)(478),
      output(27) => mem_array(27)(478),
      output(28) => mem_array(28)(478),
      output(29) => mem_array(29)(478),
      output(30) => mem_array(30)(478),
      output(31) => mem_array(31)(478),
      output(32) => mem_array(32)(478),
      output(33) => mem_array(33)(478),
      output(34) => mem_array(34)(478),
      output(35) => mem_array(35)(478)
      );
  rom479 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(479),
      output(0)  => mem_array(0)(479),
      output(1)  => mem_array(1)(479),
      output(2)  => mem_array(2)(479),
      output(3)  => mem_array(3)(479),
      output(4)  => mem_array(4)(479),
      output(5)  => mem_array(5)(479),
      output(6)  => mem_array(6)(479),
      output(7)  => mem_array(7)(479),
      output(8)  => mem_array(8)(479),
      output(9)  => mem_array(9)(479),
      output(10) => mem_array(10)(479),
      output(11) => mem_array(11)(479),
      output(12) => mem_array(12)(479),
      output(13) => mem_array(13)(479),
      output(14) => mem_array(14)(479),
      output(15) => mem_array(15)(479),
      output(16) => mem_array(16)(479),
      output(17) => mem_array(17)(479),
      output(18) => mem_array(18)(479),
      output(19) => mem_array(19)(479),
      output(20) => mem_array(20)(479),
      output(21) => mem_array(21)(479),
      output(22) => mem_array(22)(479),
      output(23) => mem_array(23)(479),
      output(24) => mem_array(24)(479),
      output(25) => mem_array(25)(479),
      output(26) => mem_array(26)(479),
      output(27) => mem_array(27)(479),
      output(28) => mem_array(28)(479),
      output(29) => mem_array(29)(479),
      output(30) => mem_array(30)(479),
      output(31) => mem_array(31)(479),
      output(32) => mem_array(32)(479),
      output(33) => mem_array(33)(479),
      output(34) => mem_array(34)(479),
      output(35) => mem_array(35)(479)
      );
  rom480 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(480),
      output(0)  => mem_array(0)(480),
      output(1)  => mem_array(1)(480),
      output(2)  => mem_array(2)(480),
      output(3)  => mem_array(3)(480),
      output(4)  => mem_array(4)(480),
      output(5)  => mem_array(5)(480),
      output(6)  => mem_array(6)(480),
      output(7)  => mem_array(7)(480),
      output(8)  => mem_array(8)(480),
      output(9)  => mem_array(9)(480),
      output(10) => mem_array(10)(480),
      output(11) => mem_array(11)(480),
      output(12) => mem_array(12)(480),
      output(13) => mem_array(13)(480),
      output(14) => mem_array(14)(480),
      output(15) => mem_array(15)(480),
      output(16) => mem_array(16)(480),
      output(17) => mem_array(17)(480),
      output(18) => mem_array(18)(480),
      output(19) => mem_array(19)(480),
      output(20) => mem_array(20)(480),
      output(21) => mem_array(21)(480),
      output(22) => mem_array(22)(480),
      output(23) => mem_array(23)(480),
      output(24) => mem_array(24)(480),
      output(25) => mem_array(25)(480),
      output(26) => mem_array(26)(480),
      output(27) => mem_array(27)(480),
      output(28) => mem_array(28)(480),
      output(29) => mem_array(29)(480),
      output(30) => mem_array(30)(480),
      output(31) => mem_array(31)(480),
      output(32) => mem_array(32)(480),
      output(33) => mem_array(33)(480),
      output(34) => mem_array(34)(480),
      output(35) => mem_array(35)(480)
      );
  rom481 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(481),
      output(0)  => mem_array(0)(481),
      output(1)  => mem_array(1)(481),
      output(2)  => mem_array(2)(481),
      output(3)  => mem_array(3)(481),
      output(4)  => mem_array(4)(481),
      output(5)  => mem_array(5)(481),
      output(6)  => mem_array(6)(481),
      output(7)  => mem_array(7)(481),
      output(8)  => mem_array(8)(481),
      output(9)  => mem_array(9)(481),
      output(10) => mem_array(10)(481),
      output(11) => mem_array(11)(481),
      output(12) => mem_array(12)(481),
      output(13) => mem_array(13)(481),
      output(14) => mem_array(14)(481),
      output(15) => mem_array(15)(481),
      output(16) => mem_array(16)(481),
      output(17) => mem_array(17)(481),
      output(18) => mem_array(18)(481),
      output(19) => mem_array(19)(481),
      output(20) => mem_array(20)(481),
      output(21) => mem_array(21)(481),
      output(22) => mem_array(22)(481),
      output(23) => mem_array(23)(481),
      output(24) => mem_array(24)(481),
      output(25) => mem_array(25)(481),
      output(26) => mem_array(26)(481),
      output(27) => mem_array(27)(481),
      output(28) => mem_array(28)(481),
      output(29) => mem_array(29)(481),
      output(30) => mem_array(30)(481),
      output(31) => mem_array(31)(481),
      output(32) => mem_array(32)(481),
      output(33) => mem_array(33)(481),
      output(34) => mem_array(34)(481),
      output(35) => mem_array(35)(481)
      );
  rom482 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(482),
      output(0)  => mem_array(0)(482),
      output(1)  => mem_array(1)(482),
      output(2)  => mem_array(2)(482),
      output(3)  => mem_array(3)(482),
      output(4)  => mem_array(4)(482),
      output(5)  => mem_array(5)(482),
      output(6)  => mem_array(6)(482),
      output(7)  => mem_array(7)(482),
      output(8)  => mem_array(8)(482),
      output(9)  => mem_array(9)(482),
      output(10) => mem_array(10)(482),
      output(11) => mem_array(11)(482),
      output(12) => mem_array(12)(482),
      output(13) => mem_array(13)(482),
      output(14) => mem_array(14)(482),
      output(15) => mem_array(15)(482),
      output(16) => mem_array(16)(482),
      output(17) => mem_array(17)(482),
      output(18) => mem_array(18)(482),
      output(19) => mem_array(19)(482),
      output(20) => mem_array(20)(482),
      output(21) => mem_array(21)(482),
      output(22) => mem_array(22)(482),
      output(23) => mem_array(23)(482),
      output(24) => mem_array(24)(482),
      output(25) => mem_array(25)(482),
      output(26) => mem_array(26)(482),
      output(27) => mem_array(27)(482),
      output(28) => mem_array(28)(482),
      output(29) => mem_array(29)(482),
      output(30) => mem_array(30)(482),
      output(31) => mem_array(31)(482),
      output(32) => mem_array(32)(482),
      output(33) => mem_array(33)(482),
      output(34) => mem_array(34)(482),
      output(35) => mem_array(35)(482)
      );
  rom483 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(483),
      output(0)  => mem_array(0)(483),
      output(1)  => mem_array(1)(483),
      output(2)  => mem_array(2)(483),
      output(3)  => mem_array(3)(483),
      output(4)  => mem_array(4)(483),
      output(5)  => mem_array(5)(483),
      output(6)  => mem_array(6)(483),
      output(7)  => mem_array(7)(483),
      output(8)  => mem_array(8)(483),
      output(9)  => mem_array(9)(483),
      output(10) => mem_array(10)(483),
      output(11) => mem_array(11)(483),
      output(12) => mem_array(12)(483),
      output(13) => mem_array(13)(483),
      output(14) => mem_array(14)(483),
      output(15) => mem_array(15)(483),
      output(16) => mem_array(16)(483),
      output(17) => mem_array(17)(483),
      output(18) => mem_array(18)(483),
      output(19) => mem_array(19)(483),
      output(20) => mem_array(20)(483),
      output(21) => mem_array(21)(483),
      output(22) => mem_array(22)(483),
      output(23) => mem_array(23)(483),
      output(24) => mem_array(24)(483),
      output(25) => mem_array(25)(483),
      output(26) => mem_array(26)(483),
      output(27) => mem_array(27)(483),
      output(28) => mem_array(28)(483),
      output(29) => mem_array(29)(483),
      output(30) => mem_array(30)(483),
      output(31) => mem_array(31)(483),
      output(32) => mem_array(32)(483),
      output(33) => mem_array(33)(483),
      output(34) => mem_array(34)(483),
      output(35) => mem_array(35)(483)
      );
  rom484 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(484),
      output(0)  => mem_array(0)(484),
      output(1)  => mem_array(1)(484),
      output(2)  => mem_array(2)(484),
      output(3)  => mem_array(3)(484),
      output(4)  => mem_array(4)(484),
      output(5)  => mem_array(5)(484),
      output(6)  => mem_array(6)(484),
      output(7)  => mem_array(7)(484),
      output(8)  => mem_array(8)(484),
      output(9)  => mem_array(9)(484),
      output(10) => mem_array(10)(484),
      output(11) => mem_array(11)(484),
      output(12) => mem_array(12)(484),
      output(13) => mem_array(13)(484),
      output(14) => mem_array(14)(484),
      output(15) => mem_array(15)(484),
      output(16) => mem_array(16)(484),
      output(17) => mem_array(17)(484),
      output(18) => mem_array(18)(484),
      output(19) => mem_array(19)(484),
      output(20) => mem_array(20)(484),
      output(21) => mem_array(21)(484),
      output(22) => mem_array(22)(484),
      output(23) => mem_array(23)(484),
      output(24) => mem_array(24)(484),
      output(25) => mem_array(25)(484),
      output(26) => mem_array(26)(484),
      output(27) => mem_array(27)(484),
      output(28) => mem_array(28)(484),
      output(29) => mem_array(29)(484),
      output(30) => mem_array(30)(484),
      output(31) => mem_array(31)(484),
      output(32) => mem_array(32)(484),
      output(33) => mem_array(33)(484),
      output(34) => mem_array(34)(484),
      output(35) => mem_array(35)(484)
      );
  rom485 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(485),
      output(0)  => mem_array(0)(485),
      output(1)  => mem_array(1)(485),
      output(2)  => mem_array(2)(485),
      output(3)  => mem_array(3)(485),
      output(4)  => mem_array(4)(485),
      output(5)  => mem_array(5)(485),
      output(6)  => mem_array(6)(485),
      output(7)  => mem_array(7)(485),
      output(8)  => mem_array(8)(485),
      output(9)  => mem_array(9)(485),
      output(10) => mem_array(10)(485),
      output(11) => mem_array(11)(485),
      output(12) => mem_array(12)(485),
      output(13) => mem_array(13)(485),
      output(14) => mem_array(14)(485),
      output(15) => mem_array(15)(485),
      output(16) => mem_array(16)(485),
      output(17) => mem_array(17)(485),
      output(18) => mem_array(18)(485),
      output(19) => mem_array(19)(485),
      output(20) => mem_array(20)(485),
      output(21) => mem_array(21)(485),
      output(22) => mem_array(22)(485),
      output(23) => mem_array(23)(485),
      output(24) => mem_array(24)(485),
      output(25) => mem_array(25)(485),
      output(26) => mem_array(26)(485),
      output(27) => mem_array(27)(485),
      output(28) => mem_array(28)(485),
      output(29) => mem_array(29)(485),
      output(30) => mem_array(30)(485),
      output(31) => mem_array(31)(485),
      output(32) => mem_array(32)(485),
      output(33) => mem_array(33)(485),
      output(34) => mem_array(34)(485),
      output(35) => mem_array(35)(485)
      );
  rom486 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(486),
      output(0)  => mem_array(0)(486),
      output(1)  => mem_array(1)(486),
      output(2)  => mem_array(2)(486),
      output(3)  => mem_array(3)(486),
      output(4)  => mem_array(4)(486),
      output(5)  => mem_array(5)(486),
      output(6)  => mem_array(6)(486),
      output(7)  => mem_array(7)(486),
      output(8)  => mem_array(8)(486),
      output(9)  => mem_array(9)(486),
      output(10) => mem_array(10)(486),
      output(11) => mem_array(11)(486),
      output(12) => mem_array(12)(486),
      output(13) => mem_array(13)(486),
      output(14) => mem_array(14)(486),
      output(15) => mem_array(15)(486),
      output(16) => mem_array(16)(486),
      output(17) => mem_array(17)(486),
      output(18) => mem_array(18)(486),
      output(19) => mem_array(19)(486),
      output(20) => mem_array(20)(486),
      output(21) => mem_array(21)(486),
      output(22) => mem_array(22)(486),
      output(23) => mem_array(23)(486),
      output(24) => mem_array(24)(486),
      output(25) => mem_array(25)(486),
      output(26) => mem_array(26)(486),
      output(27) => mem_array(27)(486),
      output(28) => mem_array(28)(486),
      output(29) => mem_array(29)(486),
      output(30) => mem_array(30)(486),
      output(31) => mem_array(31)(486),
      output(32) => mem_array(32)(486),
      output(33) => mem_array(33)(486),
      output(34) => mem_array(34)(486),
      output(35) => mem_array(35)(486)
      );
  rom487 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(487),
      output(0)  => mem_array(0)(487),
      output(1)  => mem_array(1)(487),
      output(2)  => mem_array(2)(487),
      output(3)  => mem_array(3)(487),
      output(4)  => mem_array(4)(487),
      output(5)  => mem_array(5)(487),
      output(6)  => mem_array(6)(487),
      output(7)  => mem_array(7)(487),
      output(8)  => mem_array(8)(487),
      output(9)  => mem_array(9)(487),
      output(10) => mem_array(10)(487),
      output(11) => mem_array(11)(487),
      output(12) => mem_array(12)(487),
      output(13) => mem_array(13)(487),
      output(14) => mem_array(14)(487),
      output(15) => mem_array(15)(487),
      output(16) => mem_array(16)(487),
      output(17) => mem_array(17)(487),
      output(18) => mem_array(18)(487),
      output(19) => mem_array(19)(487),
      output(20) => mem_array(20)(487),
      output(21) => mem_array(21)(487),
      output(22) => mem_array(22)(487),
      output(23) => mem_array(23)(487),
      output(24) => mem_array(24)(487),
      output(25) => mem_array(25)(487),
      output(26) => mem_array(26)(487),
      output(27) => mem_array(27)(487),
      output(28) => mem_array(28)(487),
      output(29) => mem_array(29)(487),
      output(30) => mem_array(30)(487),
      output(31) => mem_array(31)(487),
      output(32) => mem_array(32)(487),
      output(33) => mem_array(33)(487),
      output(34) => mem_array(34)(487),
      output(35) => mem_array(35)(487)
      );
  rom488 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(488),
      output(0)  => mem_array(0)(488),
      output(1)  => mem_array(1)(488),
      output(2)  => mem_array(2)(488),
      output(3)  => mem_array(3)(488),
      output(4)  => mem_array(4)(488),
      output(5)  => mem_array(5)(488),
      output(6)  => mem_array(6)(488),
      output(7)  => mem_array(7)(488),
      output(8)  => mem_array(8)(488),
      output(9)  => mem_array(9)(488),
      output(10) => mem_array(10)(488),
      output(11) => mem_array(11)(488),
      output(12) => mem_array(12)(488),
      output(13) => mem_array(13)(488),
      output(14) => mem_array(14)(488),
      output(15) => mem_array(15)(488),
      output(16) => mem_array(16)(488),
      output(17) => mem_array(17)(488),
      output(18) => mem_array(18)(488),
      output(19) => mem_array(19)(488),
      output(20) => mem_array(20)(488),
      output(21) => mem_array(21)(488),
      output(22) => mem_array(22)(488),
      output(23) => mem_array(23)(488),
      output(24) => mem_array(24)(488),
      output(25) => mem_array(25)(488),
      output(26) => mem_array(26)(488),
      output(27) => mem_array(27)(488),
      output(28) => mem_array(28)(488),
      output(29) => mem_array(29)(488),
      output(30) => mem_array(30)(488),
      output(31) => mem_array(31)(488),
      output(32) => mem_array(32)(488),
      output(33) => mem_array(33)(488),
      output(34) => mem_array(34)(488),
      output(35) => mem_array(35)(488)
      );
  rom489 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(489),
      output(0)  => mem_array(0)(489),
      output(1)  => mem_array(1)(489),
      output(2)  => mem_array(2)(489),
      output(3)  => mem_array(3)(489),
      output(4)  => mem_array(4)(489),
      output(5)  => mem_array(5)(489),
      output(6)  => mem_array(6)(489),
      output(7)  => mem_array(7)(489),
      output(8)  => mem_array(8)(489),
      output(9)  => mem_array(9)(489),
      output(10) => mem_array(10)(489),
      output(11) => mem_array(11)(489),
      output(12) => mem_array(12)(489),
      output(13) => mem_array(13)(489),
      output(14) => mem_array(14)(489),
      output(15) => mem_array(15)(489),
      output(16) => mem_array(16)(489),
      output(17) => mem_array(17)(489),
      output(18) => mem_array(18)(489),
      output(19) => mem_array(19)(489),
      output(20) => mem_array(20)(489),
      output(21) => mem_array(21)(489),
      output(22) => mem_array(22)(489),
      output(23) => mem_array(23)(489),
      output(24) => mem_array(24)(489),
      output(25) => mem_array(25)(489),
      output(26) => mem_array(26)(489),
      output(27) => mem_array(27)(489),
      output(28) => mem_array(28)(489),
      output(29) => mem_array(29)(489),
      output(30) => mem_array(30)(489),
      output(31) => mem_array(31)(489),
      output(32) => mem_array(32)(489),
      output(33) => mem_array(33)(489),
      output(34) => mem_array(34)(489),
      output(35) => mem_array(35)(489)
      );
  rom490 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(490),
      output(0)  => mem_array(0)(490),
      output(1)  => mem_array(1)(490),
      output(2)  => mem_array(2)(490),
      output(3)  => mem_array(3)(490),
      output(4)  => mem_array(4)(490),
      output(5)  => mem_array(5)(490),
      output(6)  => mem_array(6)(490),
      output(7)  => mem_array(7)(490),
      output(8)  => mem_array(8)(490),
      output(9)  => mem_array(9)(490),
      output(10) => mem_array(10)(490),
      output(11) => mem_array(11)(490),
      output(12) => mem_array(12)(490),
      output(13) => mem_array(13)(490),
      output(14) => mem_array(14)(490),
      output(15) => mem_array(15)(490),
      output(16) => mem_array(16)(490),
      output(17) => mem_array(17)(490),
      output(18) => mem_array(18)(490),
      output(19) => mem_array(19)(490),
      output(20) => mem_array(20)(490),
      output(21) => mem_array(21)(490),
      output(22) => mem_array(22)(490),
      output(23) => mem_array(23)(490),
      output(24) => mem_array(24)(490),
      output(25) => mem_array(25)(490),
      output(26) => mem_array(26)(490),
      output(27) => mem_array(27)(490),
      output(28) => mem_array(28)(490),
      output(29) => mem_array(29)(490),
      output(30) => mem_array(30)(490),
      output(31) => mem_array(31)(490),
      output(32) => mem_array(32)(490),
      output(33) => mem_array(33)(490),
      output(34) => mem_array(34)(490),
      output(35) => mem_array(35)(490)
      );
  rom491 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(491),
      output(0)  => mem_array(0)(491),
      output(1)  => mem_array(1)(491),
      output(2)  => mem_array(2)(491),
      output(3)  => mem_array(3)(491),
      output(4)  => mem_array(4)(491),
      output(5)  => mem_array(5)(491),
      output(6)  => mem_array(6)(491),
      output(7)  => mem_array(7)(491),
      output(8)  => mem_array(8)(491),
      output(9)  => mem_array(9)(491),
      output(10) => mem_array(10)(491),
      output(11) => mem_array(11)(491),
      output(12) => mem_array(12)(491),
      output(13) => mem_array(13)(491),
      output(14) => mem_array(14)(491),
      output(15) => mem_array(15)(491),
      output(16) => mem_array(16)(491),
      output(17) => mem_array(17)(491),
      output(18) => mem_array(18)(491),
      output(19) => mem_array(19)(491),
      output(20) => mem_array(20)(491),
      output(21) => mem_array(21)(491),
      output(22) => mem_array(22)(491),
      output(23) => mem_array(23)(491),
      output(24) => mem_array(24)(491),
      output(25) => mem_array(25)(491),
      output(26) => mem_array(26)(491),
      output(27) => mem_array(27)(491),
      output(28) => mem_array(28)(491),
      output(29) => mem_array(29)(491),
      output(30) => mem_array(30)(491),
      output(31) => mem_array(31)(491),
      output(32) => mem_array(32)(491),
      output(33) => mem_array(33)(491),
      output(34) => mem_array(34)(491),
      output(35) => mem_array(35)(491)
      );
  rom492 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(492),
      output(0)  => mem_array(0)(492),
      output(1)  => mem_array(1)(492),
      output(2)  => mem_array(2)(492),
      output(3)  => mem_array(3)(492),
      output(4)  => mem_array(4)(492),
      output(5)  => mem_array(5)(492),
      output(6)  => mem_array(6)(492),
      output(7)  => mem_array(7)(492),
      output(8)  => mem_array(8)(492),
      output(9)  => mem_array(9)(492),
      output(10) => mem_array(10)(492),
      output(11) => mem_array(11)(492),
      output(12) => mem_array(12)(492),
      output(13) => mem_array(13)(492),
      output(14) => mem_array(14)(492),
      output(15) => mem_array(15)(492),
      output(16) => mem_array(16)(492),
      output(17) => mem_array(17)(492),
      output(18) => mem_array(18)(492),
      output(19) => mem_array(19)(492),
      output(20) => mem_array(20)(492),
      output(21) => mem_array(21)(492),
      output(22) => mem_array(22)(492),
      output(23) => mem_array(23)(492),
      output(24) => mem_array(24)(492),
      output(25) => mem_array(25)(492),
      output(26) => mem_array(26)(492),
      output(27) => mem_array(27)(492),
      output(28) => mem_array(28)(492),
      output(29) => mem_array(29)(492),
      output(30) => mem_array(30)(492),
      output(31) => mem_array(31)(492),
      output(32) => mem_array(32)(492),
      output(33) => mem_array(33)(492),
      output(34) => mem_array(34)(492),
      output(35) => mem_array(35)(492)
      );
  rom493 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(493),
      output(0)  => mem_array(0)(493),
      output(1)  => mem_array(1)(493),
      output(2)  => mem_array(2)(493),
      output(3)  => mem_array(3)(493),
      output(4)  => mem_array(4)(493),
      output(5)  => mem_array(5)(493),
      output(6)  => mem_array(6)(493),
      output(7)  => mem_array(7)(493),
      output(8)  => mem_array(8)(493),
      output(9)  => mem_array(9)(493),
      output(10) => mem_array(10)(493),
      output(11) => mem_array(11)(493),
      output(12) => mem_array(12)(493),
      output(13) => mem_array(13)(493),
      output(14) => mem_array(14)(493),
      output(15) => mem_array(15)(493),
      output(16) => mem_array(16)(493),
      output(17) => mem_array(17)(493),
      output(18) => mem_array(18)(493),
      output(19) => mem_array(19)(493),
      output(20) => mem_array(20)(493),
      output(21) => mem_array(21)(493),
      output(22) => mem_array(22)(493),
      output(23) => mem_array(23)(493),
      output(24) => mem_array(24)(493),
      output(25) => mem_array(25)(493),
      output(26) => mem_array(26)(493),
      output(27) => mem_array(27)(493),
      output(28) => mem_array(28)(493),
      output(29) => mem_array(29)(493),
      output(30) => mem_array(30)(493),
      output(31) => mem_array(31)(493),
      output(32) => mem_array(32)(493),
      output(33) => mem_array(33)(493),
      output(34) => mem_array(34)(493),
      output(35) => mem_array(35)(493)
      );
  rom494 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(494),
      output(0)  => mem_array(0)(494),
      output(1)  => mem_array(1)(494),
      output(2)  => mem_array(2)(494),
      output(3)  => mem_array(3)(494),
      output(4)  => mem_array(4)(494),
      output(5)  => mem_array(5)(494),
      output(6)  => mem_array(6)(494),
      output(7)  => mem_array(7)(494),
      output(8)  => mem_array(8)(494),
      output(9)  => mem_array(9)(494),
      output(10) => mem_array(10)(494),
      output(11) => mem_array(11)(494),
      output(12) => mem_array(12)(494),
      output(13) => mem_array(13)(494),
      output(14) => mem_array(14)(494),
      output(15) => mem_array(15)(494),
      output(16) => mem_array(16)(494),
      output(17) => mem_array(17)(494),
      output(18) => mem_array(18)(494),
      output(19) => mem_array(19)(494),
      output(20) => mem_array(20)(494),
      output(21) => mem_array(21)(494),
      output(22) => mem_array(22)(494),
      output(23) => mem_array(23)(494),
      output(24) => mem_array(24)(494),
      output(25) => mem_array(25)(494),
      output(26) => mem_array(26)(494),
      output(27) => mem_array(27)(494),
      output(28) => mem_array(28)(494),
      output(29) => mem_array(29)(494),
      output(30) => mem_array(30)(494),
      output(31) => mem_array(31)(494),
      output(32) => mem_array(32)(494),
      output(33) => mem_array(33)(494),
      output(34) => mem_array(34)(494),
      output(35) => mem_array(35)(494)
      );
  rom495 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(495),
      output(0)  => mem_array(0)(495),
      output(1)  => mem_array(1)(495),
      output(2)  => mem_array(2)(495),
      output(3)  => mem_array(3)(495),
      output(4)  => mem_array(4)(495),
      output(5)  => mem_array(5)(495),
      output(6)  => mem_array(6)(495),
      output(7)  => mem_array(7)(495),
      output(8)  => mem_array(8)(495),
      output(9)  => mem_array(9)(495),
      output(10) => mem_array(10)(495),
      output(11) => mem_array(11)(495),
      output(12) => mem_array(12)(495),
      output(13) => mem_array(13)(495),
      output(14) => mem_array(14)(495),
      output(15) => mem_array(15)(495),
      output(16) => mem_array(16)(495),
      output(17) => mem_array(17)(495),
      output(18) => mem_array(18)(495),
      output(19) => mem_array(19)(495),
      output(20) => mem_array(20)(495),
      output(21) => mem_array(21)(495),
      output(22) => mem_array(22)(495),
      output(23) => mem_array(23)(495),
      output(24) => mem_array(24)(495),
      output(25) => mem_array(25)(495),
      output(26) => mem_array(26)(495),
      output(27) => mem_array(27)(495),
      output(28) => mem_array(28)(495),
      output(29) => mem_array(29)(495),
      output(30) => mem_array(30)(495),
      output(31) => mem_array(31)(495),
      output(32) => mem_array(32)(495),
      output(33) => mem_array(33)(495),
      output(34) => mem_array(34)(495),
      output(35) => mem_array(35)(495)
      );
  rom496 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(496),
      output(0)  => mem_array(0)(496),
      output(1)  => mem_array(1)(496),
      output(2)  => mem_array(2)(496),
      output(3)  => mem_array(3)(496),
      output(4)  => mem_array(4)(496),
      output(5)  => mem_array(5)(496),
      output(6)  => mem_array(6)(496),
      output(7)  => mem_array(7)(496),
      output(8)  => mem_array(8)(496),
      output(9)  => mem_array(9)(496),
      output(10) => mem_array(10)(496),
      output(11) => mem_array(11)(496),
      output(12) => mem_array(12)(496),
      output(13) => mem_array(13)(496),
      output(14) => mem_array(14)(496),
      output(15) => mem_array(15)(496),
      output(16) => mem_array(16)(496),
      output(17) => mem_array(17)(496),
      output(18) => mem_array(18)(496),
      output(19) => mem_array(19)(496),
      output(20) => mem_array(20)(496),
      output(21) => mem_array(21)(496),
      output(22) => mem_array(22)(496),
      output(23) => mem_array(23)(496),
      output(24) => mem_array(24)(496),
      output(25) => mem_array(25)(496),
      output(26) => mem_array(26)(496),
      output(27) => mem_array(27)(496),
      output(28) => mem_array(28)(496),
      output(29) => mem_array(29)(496),
      output(30) => mem_array(30)(496),
      output(31) => mem_array(31)(496),
      output(32) => mem_array(32)(496),
      output(33) => mem_array(33)(496),
      output(34) => mem_array(34)(496),
      output(35) => mem_array(35)(496)
      );
  rom497 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(497),
      output(0)  => mem_array(0)(497),
      output(1)  => mem_array(1)(497),
      output(2)  => mem_array(2)(497),
      output(3)  => mem_array(3)(497),
      output(4)  => mem_array(4)(497),
      output(5)  => mem_array(5)(497),
      output(6)  => mem_array(6)(497),
      output(7)  => mem_array(7)(497),
      output(8)  => mem_array(8)(497),
      output(9)  => mem_array(9)(497),
      output(10) => mem_array(10)(497),
      output(11) => mem_array(11)(497),
      output(12) => mem_array(12)(497),
      output(13) => mem_array(13)(497),
      output(14) => mem_array(14)(497),
      output(15) => mem_array(15)(497),
      output(16) => mem_array(16)(497),
      output(17) => mem_array(17)(497),
      output(18) => mem_array(18)(497),
      output(19) => mem_array(19)(497),
      output(20) => mem_array(20)(497),
      output(21) => mem_array(21)(497),
      output(22) => mem_array(22)(497),
      output(23) => mem_array(23)(497),
      output(24) => mem_array(24)(497),
      output(25) => mem_array(25)(497),
      output(26) => mem_array(26)(497),
      output(27) => mem_array(27)(497),
      output(28) => mem_array(28)(497),
      output(29) => mem_array(29)(497),
      output(30) => mem_array(30)(497),
      output(31) => mem_array(31)(497),
      output(32) => mem_array(32)(497),
      output(33) => mem_array(33)(497),
      output(34) => mem_array(34)(497),
      output(35) => mem_array(35)(497)
      );
  rom498 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(498),
      output(0)  => mem_array(0)(498),
      output(1)  => mem_array(1)(498),
      output(2)  => mem_array(2)(498),
      output(3)  => mem_array(3)(498),
      output(4)  => mem_array(4)(498),
      output(5)  => mem_array(5)(498),
      output(6)  => mem_array(6)(498),
      output(7)  => mem_array(7)(498),
      output(8)  => mem_array(8)(498),
      output(9)  => mem_array(9)(498),
      output(10) => mem_array(10)(498),
      output(11) => mem_array(11)(498),
      output(12) => mem_array(12)(498),
      output(13) => mem_array(13)(498),
      output(14) => mem_array(14)(498),
      output(15) => mem_array(15)(498),
      output(16) => mem_array(16)(498),
      output(17) => mem_array(17)(498),
      output(18) => mem_array(18)(498),
      output(19) => mem_array(19)(498),
      output(20) => mem_array(20)(498),
      output(21) => mem_array(21)(498),
      output(22) => mem_array(22)(498),
      output(23) => mem_array(23)(498),
      output(24) => mem_array(24)(498),
      output(25) => mem_array(25)(498),
      output(26) => mem_array(26)(498),
      output(27) => mem_array(27)(498),
      output(28) => mem_array(28)(498),
      output(29) => mem_array(29)(498),
      output(30) => mem_array(30)(498),
      output(31) => mem_array(31)(498),
      output(32) => mem_array(32)(498),
      output(33) => mem_array(33)(498),
      output(34) => mem_array(34)(498),
      output(35) => mem_array(35)(498)
      );
  rom499 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(499),
      output(0)  => mem_array(0)(499),
      output(1)  => mem_array(1)(499),
      output(2)  => mem_array(2)(499),
      output(3)  => mem_array(3)(499),
      output(4)  => mem_array(4)(499),
      output(5)  => mem_array(5)(499),
      output(6)  => mem_array(6)(499),
      output(7)  => mem_array(7)(499),
      output(8)  => mem_array(8)(499),
      output(9)  => mem_array(9)(499),
      output(10) => mem_array(10)(499),
      output(11) => mem_array(11)(499),
      output(12) => mem_array(12)(499),
      output(13) => mem_array(13)(499),
      output(14) => mem_array(14)(499),
      output(15) => mem_array(15)(499),
      output(16) => mem_array(16)(499),
      output(17) => mem_array(17)(499),
      output(18) => mem_array(18)(499),
      output(19) => mem_array(19)(499),
      output(20) => mem_array(20)(499),
      output(21) => mem_array(21)(499),
      output(22) => mem_array(22)(499),
      output(23) => mem_array(23)(499),
      output(24) => mem_array(24)(499),
      output(25) => mem_array(25)(499),
      output(26) => mem_array(26)(499),
      output(27) => mem_array(27)(499),
      output(28) => mem_array(28)(499),
      output(29) => mem_array(29)(499),
      output(30) => mem_array(30)(499),
      output(31) => mem_array(31)(499),
      output(32) => mem_array(32)(499),
      output(33) => mem_array(33)(499),
      output(34) => mem_array(34)(499),
      output(35) => mem_array(35)(499)
      );
  rom500 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(500),
      output(0)  => mem_array(0)(500),
      output(1)  => mem_array(1)(500),
      output(2)  => mem_array(2)(500),
      output(3)  => mem_array(3)(500),
      output(4)  => mem_array(4)(500),
      output(5)  => mem_array(5)(500),
      output(6)  => mem_array(6)(500),
      output(7)  => mem_array(7)(500),
      output(8)  => mem_array(8)(500),
      output(9)  => mem_array(9)(500),
      output(10) => mem_array(10)(500),
      output(11) => mem_array(11)(500),
      output(12) => mem_array(12)(500),
      output(13) => mem_array(13)(500),
      output(14) => mem_array(14)(500),
      output(15) => mem_array(15)(500),
      output(16) => mem_array(16)(500),
      output(17) => mem_array(17)(500),
      output(18) => mem_array(18)(500),
      output(19) => mem_array(19)(500),
      output(20) => mem_array(20)(500),
      output(21) => mem_array(21)(500),
      output(22) => mem_array(22)(500),
      output(23) => mem_array(23)(500),
      output(24) => mem_array(24)(500),
      output(25) => mem_array(25)(500),
      output(26) => mem_array(26)(500),
      output(27) => mem_array(27)(500),
      output(28) => mem_array(28)(500),
      output(29) => mem_array(29)(500),
      output(30) => mem_array(30)(500),
      output(31) => mem_array(31)(500),
      output(32) => mem_array(32)(500),
      output(33) => mem_array(33)(500),
      output(34) => mem_array(34)(500),
      output(35) => mem_array(35)(500)
      );
  rom501 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(501),
      output(0)  => mem_array(0)(501),
      output(1)  => mem_array(1)(501),
      output(2)  => mem_array(2)(501),
      output(3)  => mem_array(3)(501),
      output(4)  => mem_array(4)(501),
      output(5)  => mem_array(5)(501),
      output(6)  => mem_array(6)(501),
      output(7)  => mem_array(7)(501),
      output(8)  => mem_array(8)(501),
      output(9)  => mem_array(9)(501),
      output(10) => mem_array(10)(501),
      output(11) => mem_array(11)(501),
      output(12) => mem_array(12)(501),
      output(13) => mem_array(13)(501),
      output(14) => mem_array(14)(501),
      output(15) => mem_array(15)(501),
      output(16) => mem_array(16)(501),
      output(17) => mem_array(17)(501),
      output(18) => mem_array(18)(501),
      output(19) => mem_array(19)(501),
      output(20) => mem_array(20)(501),
      output(21) => mem_array(21)(501),
      output(22) => mem_array(22)(501),
      output(23) => mem_array(23)(501),
      output(24) => mem_array(24)(501),
      output(25) => mem_array(25)(501),
      output(26) => mem_array(26)(501),
      output(27) => mem_array(27)(501),
      output(28) => mem_array(28)(501),
      output(29) => mem_array(29)(501),
      output(30) => mem_array(30)(501),
      output(31) => mem_array(31)(501),
      output(32) => mem_array(32)(501),
      output(33) => mem_array(33)(501),
      output(34) => mem_array(34)(501),
      output(35) => mem_array(35)(501)
      );
  rom502 : entity work.rom
    generic map (
      bits  => 36,
      value => "011111110000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(502),
      output(0)  => mem_array(0)(502),
      output(1)  => mem_array(1)(502),
      output(2)  => mem_array(2)(502),
      output(3)  => mem_array(3)(502),
      output(4)  => mem_array(4)(502),
      output(5)  => mem_array(5)(502),
      output(6)  => mem_array(6)(502),
      output(7)  => mem_array(7)(502),
      output(8)  => mem_array(8)(502),
      output(9)  => mem_array(9)(502),
      output(10) => mem_array(10)(502),
      output(11) => mem_array(11)(502),
      output(12) => mem_array(12)(502),
      output(13) => mem_array(13)(502),
      output(14) => mem_array(14)(502),
      output(15) => mem_array(15)(502),
      output(16) => mem_array(16)(502),
      output(17) => mem_array(17)(502),
      output(18) => mem_array(18)(502),
      output(19) => mem_array(19)(502),
      output(20) => mem_array(20)(502),
      output(21) => mem_array(21)(502),
      output(22) => mem_array(22)(502),
      output(23) => mem_array(23)(502),
      output(24) => mem_array(24)(502),
      output(25) => mem_array(25)(502),
      output(26) => mem_array(26)(502),
      output(27) => mem_array(27)(502),
      output(28) => mem_array(28)(502),
      output(29) => mem_array(29)(502),
      output(30) => mem_array(30)(502),
      output(31) => mem_array(31)(502),
      output(32) => mem_array(32)(502),
      output(33) => mem_array(33)(502),
      output(34) => mem_array(34)(502),
      output(35) => mem_array(35)(502)
      );
  rom503 : entity work.rom
    generic map (
      bits  => 36,
      value => "000001111111000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(503),
      output(0)  => mem_array(0)(503),
      output(1)  => mem_array(1)(503),
      output(2)  => mem_array(2)(503),
      output(3)  => mem_array(3)(503),
      output(4)  => mem_array(4)(503),
      output(5)  => mem_array(5)(503),
      output(6)  => mem_array(6)(503),
      output(7)  => mem_array(7)(503),
      output(8)  => mem_array(8)(503),
      output(9)  => mem_array(9)(503),
      output(10) => mem_array(10)(503),
      output(11) => mem_array(11)(503),
      output(12) => mem_array(12)(503),
      output(13) => mem_array(13)(503),
      output(14) => mem_array(14)(503),
      output(15) => mem_array(15)(503),
      output(16) => mem_array(16)(503),
      output(17) => mem_array(17)(503),
      output(18) => mem_array(18)(503),
      output(19) => mem_array(19)(503),
      output(20) => mem_array(20)(503),
      output(21) => mem_array(21)(503),
      output(22) => mem_array(22)(503),
      output(23) => mem_array(23)(503),
      output(24) => mem_array(24)(503),
      output(25) => mem_array(25)(503),
      output(26) => mem_array(26)(503),
      output(27) => mem_array(27)(503),
      output(28) => mem_array(28)(503),
      output(29) => mem_array(29)(503),
      output(30) => mem_array(30)(503),
      output(31) => mem_array(31)(503),
      output(32) => mem_array(32)(503),
      output(33) => mem_array(33)(503),
      output(34) => mem_array(34)(503),
      output(35) => mem_array(35)(503)
      );
  rom504 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000111111100000000000000000000")
    port map (
      enable_o   => mem_enable_lines(504),
      output(0)  => mem_array(0)(504),
      output(1)  => mem_array(1)(504),
      output(2)  => mem_array(2)(504),
      output(3)  => mem_array(3)(504),
      output(4)  => mem_array(4)(504),
      output(5)  => mem_array(5)(504),
      output(6)  => mem_array(6)(504),
      output(7)  => mem_array(7)(504),
      output(8)  => mem_array(8)(504),
      output(9)  => mem_array(9)(504),
      output(10) => mem_array(10)(504),
      output(11) => mem_array(11)(504),
      output(12) => mem_array(12)(504),
      output(13) => mem_array(13)(504),
      output(14) => mem_array(14)(504),
      output(15) => mem_array(15)(504),
      output(16) => mem_array(16)(504),
      output(17) => mem_array(17)(504),
      output(18) => mem_array(18)(504),
      output(19) => mem_array(19)(504),
      output(20) => mem_array(20)(504),
      output(21) => mem_array(21)(504),
      output(22) => mem_array(22)(504),
      output(23) => mem_array(23)(504),
      output(24) => mem_array(24)(504),
      output(25) => mem_array(25)(504),
      output(26) => mem_array(26)(504),
      output(27) => mem_array(27)(504),
      output(28) => mem_array(28)(504),
      output(29) => mem_array(29)(504),
      output(30) => mem_array(30)(504),
      output(31) => mem_array(31)(504),
      output(32) => mem_array(32)(504),
      output(33) => mem_array(33)(504),
      output(34) => mem_array(34)(504),
      output(35) => mem_array(35)(504)
      );
  rom505 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000011111110000000000000000")
    port map (
      enable_o   => mem_enable_lines(505),
      output(0)  => mem_array(0)(505),
      output(1)  => mem_array(1)(505),
      output(2)  => mem_array(2)(505),
      output(3)  => mem_array(3)(505),
      output(4)  => mem_array(4)(505),
      output(5)  => mem_array(5)(505),
      output(6)  => mem_array(6)(505),
      output(7)  => mem_array(7)(505),
      output(8)  => mem_array(8)(505),
      output(9)  => mem_array(9)(505),
      output(10) => mem_array(10)(505),
      output(11) => mem_array(11)(505),
      output(12) => mem_array(12)(505),
      output(13) => mem_array(13)(505),
      output(14) => mem_array(14)(505),
      output(15) => mem_array(15)(505),
      output(16) => mem_array(16)(505),
      output(17) => mem_array(17)(505),
      output(18) => mem_array(18)(505),
      output(19) => mem_array(19)(505),
      output(20) => mem_array(20)(505),
      output(21) => mem_array(21)(505),
      output(22) => mem_array(22)(505),
      output(23) => mem_array(23)(505),
      output(24) => mem_array(24)(505),
      output(25) => mem_array(25)(505),
      output(26) => mem_array(26)(505),
      output(27) => mem_array(27)(505),
      output(28) => mem_array(28)(505),
      output(29) => mem_array(29)(505),
      output(30) => mem_array(30)(505),
      output(31) => mem_array(31)(505),
      output(32) => mem_array(32)(505),
      output(33) => mem_array(33)(505),
      output(34) => mem_array(34)(505),
      output(35) => mem_array(35)(505)
      );
  rom506 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000001111111000000000000")
    port map (
      enable_o   => mem_enable_lines(506),
      output(0)  => mem_array(0)(506),
      output(1)  => mem_array(1)(506),
      output(2)  => mem_array(2)(506),
      output(3)  => mem_array(3)(506),
      output(4)  => mem_array(4)(506),
      output(5)  => mem_array(5)(506),
      output(6)  => mem_array(6)(506),
      output(7)  => mem_array(7)(506),
      output(8)  => mem_array(8)(506),
      output(9)  => mem_array(9)(506),
      output(10) => mem_array(10)(506),
      output(11) => mem_array(11)(506),
      output(12) => mem_array(12)(506),
      output(13) => mem_array(13)(506),
      output(14) => mem_array(14)(506),
      output(15) => mem_array(15)(506),
      output(16) => mem_array(16)(506),
      output(17) => mem_array(17)(506),
      output(18) => mem_array(18)(506),
      output(19) => mem_array(19)(506),
      output(20) => mem_array(20)(506),
      output(21) => mem_array(21)(506),
      output(22) => mem_array(22)(506),
      output(23) => mem_array(23)(506),
      output(24) => mem_array(24)(506),
      output(25) => mem_array(25)(506),
      output(26) => mem_array(26)(506),
      output(27) => mem_array(27)(506),
      output(28) => mem_array(28)(506),
      output(29) => mem_array(29)(506),
      output(30) => mem_array(30)(506),
      output(31) => mem_array(31)(506),
      output(32) => mem_array(32)(506),
      output(33) => mem_array(33)(506),
      output(34) => mem_array(34)(506),
      output(35) => mem_array(35)(506)
      );
  rom507 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000111111100000000")
    port map (
      enable_o   => mem_enable_lines(507),
      output(0)  => mem_array(0)(507),
      output(1)  => mem_array(1)(507),
      output(2)  => mem_array(2)(507),
      output(3)  => mem_array(3)(507),
      output(4)  => mem_array(4)(507),
      output(5)  => mem_array(5)(507),
      output(6)  => mem_array(6)(507),
      output(7)  => mem_array(7)(507),
      output(8)  => mem_array(8)(507),
      output(9)  => mem_array(9)(507),
      output(10) => mem_array(10)(507),
      output(11) => mem_array(11)(507),
      output(12) => mem_array(12)(507),
      output(13) => mem_array(13)(507),
      output(14) => mem_array(14)(507),
      output(15) => mem_array(15)(507),
      output(16) => mem_array(16)(507),
      output(17) => mem_array(17)(507),
      output(18) => mem_array(18)(507),
      output(19) => mem_array(19)(507),
      output(20) => mem_array(20)(507),
      output(21) => mem_array(21)(507),
      output(22) => mem_array(22)(507),
      output(23) => mem_array(23)(507),
      output(24) => mem_array(24)(507),
      output(25) => mem_array(25)(507),
      output(26) => mem_array(26)(507),
      output(27) => mem_array(27)(507),
      output(28) => mem_array(28)(507),
      output(29) => mem_array(29)(507),
      output(30) => mem_array(30)(507),
      output(31) => mem_array(31)(507),
      output(32) => mem_array(32)(507),
      output(33) => mem_array(33)(507),
      output(34) => mem_array(34)(507),
      output(35) => mem_array(35)(507)
      );
  rom508 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000011111110000")
    port map (
      enable_o   => mem_enable_lines(508),
      output(0)  => mem_array(0)(508),
      output(1)  => mem_array(1)(508),
      output(2)  => mem_array(2)(508),
      output(3)  => mem_array(3)(508),
      output(4)  => mem_array(4)(508),
      output(5)  => mem_array(5)(508),
      output(6)  => mem_array(6)(508),
      output(7)  => mem_array(7)(508),
      output(8)  => mem_array(8)(508),
      output(9)  => mem_array(9)(508),
      output(10) => mem_array(10)(508),
      output(11) => mem_array(11)(508),
      output(12) => mem_array(12)(508),
      output(13) => mem_array(13)(508),
      output(14) => mem_array(14)(508),
      output(15) => mem_array(15)(508),
      output(16) => mem_array(16)(508),
      output(17) => mem_array(17)(508),
      output(18) => mem_array(18)(508),
      output(19) => mem_array(19)(508),
      output(20) => mem_array(20)(508),
      output(21) => mem_array(21)(508),
      output(22) => mem_array(22)(508),
      output(23) => mem_array(23)(508),
      output(24) => mem_array(24)(508),
      output(25) => mem_array(25)(508),
      output(26) => mem_array(26)(508),
      output(27) => mem_array(27)(508),
      output(28) => mem_array(28)(508),
      output(29) => mem_array(29)(508),
      output(30) => mem_array(30)(508),
      output(31) => mem_array(31)(508),
      output(32) => mem_array(32)(508),
      output(33) => mem_array(33)(508),
      output(34) => mem_array(34)(508),
      output(35) => mem_array(35)(508)
      );
  rom509 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000001111111")
    port map (
      enable_o   => mem_enable_lines(509),
      output(0)  => mem_array(0)(509),
      output(1)  => mem_array(1)(509),
      output(2)  => mem_array(2)(509),
      output(3)  => mem_array(3)(509),
      output(4)  => mem_array(4)(509),
      output(5)  => mem_array(5)(509),
      output(6)  => mem_array(6)(509),
      output(7)  => mem_array(7)(509),
      output(8)  => mem_array(8)(509),
      output(9)  => mem_array(9)(509),
      output(10) => mem_array(10)(509),
      output(11) => mem_array(11)(509),
      output(12) => mem_array(12)(509),
      output(13) => mem_array(13)(509),
      output(14) => mem_array(14)(509),
      output(15) => mem_array(15)(509),
      output(16) => mem_array(16)(509),
      output(17) => mem_array(17)(509),
      output(18) => mem_array(18)(509),
      output(19) => mem_array(19)(509),
      output(20) => mem_array(20)(509),
      output(21) => mem_array(21)(509),
      output(22) => mem_array(22)(509),
      output(23) => mem_array(23)(509),
      output(24) => mem_array(24)(509),
      output(25) => mem_array(25)(509),
      output(26) => mem_array(26)(509),
      output(27) => mem_array(27)(509),
      output(28) => mem_array(28)(509),
      output(29) => mem_array(29)(509),
      output(30) => mem_array(30)(509),
      output(31) => mem_array(31)(509),
      output(32) => mem_array(32)(509),
      output(33) => mem_array(33)(509),
      output(34) => mem_array(34)(509),
      output(35) => mem_array(35)(509)
      );
  rom510 : entity work.rom
    generic map (
      bits  => 36,
      value => "000000000000000000000000000000000111")
    port map (
      enable_o   => mem_enable_lines(510),
      output(0)  => mem_array(0)(510),
      output(1)  => mem_array(1)(510),
      output(2)  => mem_array(2)(510),
      output(3)  => mem_array(3)(510),
      output(4)  => mem_array(4)(510),
      output(5)  => mem_array(5)(510),
      output(6)  => mem_array(6)(510),
      output(7)  => mem_array(7)(510),
      output(8)  => mem_array(8)(510),
      output(9)  => mem_array(9)(510),
      output(10) => mem_array(10)(510),
      output(11) => mem_array(11)(510),
      output(12) => mem_array(12)(510),
      output(13) => mem_array(13)(510),
      output(14) => mem_array(14)(510),
      output(15) => mem_array(15)(510),
      output(16) => mem_array(16)(510),
      output(17) => mem_array(17)(510),
      output(18) => mem_array(18)(510),
      output(19) => mem_array(19)(510),
      output(20) => mem_array(20)(510),
      output(21) => mem_array(21)(510),
      output(22) => mem_array(22)(510),
      output(23) => mem_array(23)(510),
      output(24) => mem_array(24)(510),
      output(25) => mem_array(25)(510),
      output(26) => mem_array(26)(510),
      output(27) => mem_array(27)(510),
      output(28) => mem_array(28)(510),
      output(29) => mem_array(29)(510),
      output(30) => mem_array(30)(510),
      output(31) => mem_array(31)(510),
      output(32) => mem_array(32)(510),
      output(33) => mem_array(33)(510),
      output(34) => mem_array(34)(510),
      output(35) => mem_array(35)(510)
      );
  rom511 : entity work.rom
    generic map (
      bits  => 36,
      value => "111100000000000000000000000000000000")
    port map (
      enable_o   => mem_enable_lines(511),
      output(0)  => mem_array(0)(511),
      output(1)  => mem_array(1)(511),
      output(2)  => mem_array(2)(511),
      output(3)  => mem_array(3)(511),
      output(4)  => mem_array(4)(511),
      output(5)  => mem_array(5)(511),
      output(6)  => mem_array(6)(511),
      output(7)  => mem_array(7)(511),
      output(8)  => mem_array(8)(511),
      output(9)  => mem_array(9)(511),
      output(10) => mem_array(10)(511),
      output(11) => mem_array(11)(511),
      output(12) => mem_array(12)(511),
      output(13) => mem_array(13)(511),
      output(14) => mem_array(14)(511),
      output(15) => mem_array(15)(511),
      output(16) => mem_array(16)(511),
      output(17) => mem_array(17)(511),
      output(18) => mem_array(18)(511),
      output(19) => mem_array(19)(511),
      output(20) => mem_array(20)(511),
      output(21) => mem_array(21)(511),
      output(22) => mem_array(22)(511),
      output(23) => mem_array(23)(511),
      output(24) => mem_array(24)(511),
      output(25) => mem_array(25)(511),
      output(26) => mem_array(26)(511),
      output(27) => mem_array(27)(511),
      output(28) => mem_array(28)(511),
      output(29) => mem_array(29)(511),
      output(30) => mem_array(30)(511),
      output(31) => mem_array(31)(511),
      output(32) => mem_array(32)(511),
      output(33) => mem_array(33)(511),
      output(34) => mem_array(34)(511),
      output(35) => mem_array(35)(511)
      );


  -- gen: for i in 511 downto 0 generate
  --   temp_instruction <= temp_instruction or mem_array(i);
  --   test <= temp_instruction;
  -- end generate gen;
  -- instruction <= temp_instruction;

  -- gen: for i in 511 downto 0 generate
  --   temp_instruction(i) 
  -- end generate gen;

  lf : for i in 35 downto 0 generate
    instruction(i) <= or_reduce(mem_array(i));
  end generate lf;


end architecture control_store_ar;
